magic
tech scmos
timestamp 1699956227
<< nwell >>
rect 3 -173 111 -155
rect 158 -172 266 -154
rect -103 -324 -49 -306
rect -42 -324 -11 -306
rect 37 -323 91 -305
rect 98 -323 129 -305
rect 182 -322 236 -304
rect 243 -322 274 -304
rect 343 -325 443 -307
<< ntransistor >>
rect 18 -220 21 -216
rect 41 -220 44 -216
rect 72 -220 75 -216
rect 95 -220 98 -216
rect 173 -219 176 -215
rect 196 -219 199 -215
rect 227 -219 230 -215
rect 250 -219 253 -215
rect 358 -347 361 -342
rect 381 -347 384 -342
rect 404 -347 407 -342
rect 427 -347 430 -342
rect -88 -354 -85 -349
rect -65 -354 -62 -349
rect -27 -354 -24 -349
rect 52 -353 55 -348
rect 75 -353 78 -348
rect 113 -353 116 -348
rect 197 -352 200 -347
rect 220 -352 223 -347
rect 258 -352 261 -347
<< ptransistor >>
rect 18 -167 21 -161
rect 41 -167 44 -161
rect 72 -167 75 -161
rect 95 -167 98 -161
rect 173 -166 176 -160
rect 196 -166 199 -160
rect 227 -166 230 -160
rect 250 -166 253 -160
rect -88 -318 -85 -312
rect -65 -318 -62 -312
rect -27 -318 -24 -312
rect 52 -317 55 -311
rect 75 -317 78 -311
rect 113 -317 116 -311
rect 197 -316 200 -310
rect 220 -316 223 -310
rect 258 -316 261 -310
rect 358 -319 361 -313
rect 381 -319 384 -313
rect 404 -319 407 -313
rect 427 -319 430 -313
<< ndiffusion >>
rect 15 -220 18 -216
rect 21 -220 24 -216
rect 38 -220 41 -216
rect 44 -220 47 -216
rect 68 -220 72 -216
rect 75 -220 78 -216
rect 91 -220 95 -216
rect 98 -220 101 -216
rect 170 -219 173 -215
rect 176 -219 179 -215
rect 193 -219 196 -215
rect 199 -219 202 -215
rect 223 -219 227 -215
rect 230 -219 233 -215
rect 246 -219 250 -215
rect 253 -219 256 -215
rect 354 -347 358 -342
rect 361 -347 364 -342
rect 377 -347 381 -342
rect 384 -347 387 -342
rect 400 -347 404 -342
rect 407 -347 410 -342
rect 423 -347 427 -342
rect 430 -347 433 -342
rect -92 -354 -88 -349
rect -85 -354 -82 -349
rect -69 -354 -65 -349
rect -62 -354 -59 -349
rect -31 -354 -27 -349
rect -24 -354 -21 -349
rect 48 -353 52 -348
rect 55 -353 58 -348
rect 71 -353 75 -348
rect 78 -353 81 -348
rect 109 -353 113 -348
rect 116 -353 119 -348
rect 193 -352 197 -347
rect 200 -352 203 -347
rect 216 -352 220 -347
rect 223 -352 226 -347
rect 254 -352 258 -347
rect 261 -352 264 -347
<< pdiffusion >>
rect 15 -167 18 -161
rect 21 -167 24 -161
rect 38 -167 41 -161
rect 44 -167 47 -161
rect 69 -167 72 -161
rect 75 -167 78 -161
rect 92 -167 95 -161
rect 98 -167 101 -161
rect 170 -166 173 -160
rect 176 -166 179 -160
rect 193 -166 196 -160
rect 199 -166 202 -160
rect 224 -166 227 -160
rect 230 -166 233 -160
rect 247 -166 250 -160
rect 253 -166 256 -160
rect -91 -318 -88 -312
rect -85 -318 -82 -312
rect -68 -318 -65 -312
rect -62 -318 -59 -312
rect -30 -318 -27 -312
rect -24 -318 -21 -312
rect 49 -317 52 -311
rect 55 -317 58 -311
rect 72 -317 75 -311
rect 78 -317 81 -311
rect 110 -317 113 -311
rect 116 -317 119 -311
rect 194 -316 197 -310
rect 200 -316 203 -310
rect 217 -316 220 -310
rect 223 -316 226 -310
rect 255 -316 258 -310
rect 261 -316 264 -310
rect 355 -319 358 -313
rect 361 -319 364 -313
rect 378 -319 381 -313
rect 384 -319 387 -313
rect 401 -319 404 -313
rect 407 -319 410 -313
rect 424 -319 427 -313
rect 430 -319 433 -313
<< ndcontact >>
rect 10 -220 15 -216
rect 24 -220 28 -216
rect 33 -220 38 -216
rect 47 -220 51 -216
rect 64 -220 68 -216
rect 78 -220 82 -216
rect 87 -220 91 -216
rect 101 -220 105 -216
rect 165 -219 170 -215
rect 179 -219 183 -215
rect 188 -219 193 -215
rect 202 -219 206 -215
rect 219 -219 223 -215
rect 233 -219 237 -215
rect 242 -219 246 -215
rect 256 -219 260 -215
rect 350 -347 354 -342
rect 364 -347 368 -342
rect 373 -347 377 -342
rect 387 -347 391 -342
rect 396 -347 400 -342
rect 410 -347 414 -342
rect 419 -347 423 -342
rect 433 -347 437 -342
rect -96 -354 -92 -349
rect -82 -354 -78 -349
rect -73 -354 -69 -349
rect -59 -354 -55 -349
rect -35 -354 -31 -349
rect -21 -354 -17 -349
rect 44 -353 48 -348
rect 58 -353 62 -348
rect 67 -353 71 -348
rect 81 -353 85 -348
rect 105 -353 109 -348
rect 119 -353 123 -348
rect 189 -352 193 -347
rect 203 -352 207 -347
rect 212 -352 216 -347
rect 226 -352 230 -347
rect 250 -352 254 -347
rect 264 -352 268 -347
<< pdcontact >>
rect 10 -167 15 -161
rect 24 -167 28 -161
rect 33 -167 38 -161
rect 47 -167 51 -161
rect 64 -167 69 -161
rect 78 -167 82 -161
rect 87 -167 92 -161
rect 101 -167 105 -161
rect 165 -166 170 -160
rect 179 -166 183 -160
rect 188 -166 193 -160
rect 202 -166 206 -160
rect 219 -166 224 -160
rect 233 -166 237 -160
rect 242 -166 247 -160
rect 256 -166 260 -160
rect -96 -318 -91 -312
rect -82 -318 -78 -312
rect -73 -318 -68 -312
rect -59 -318 -55 -312
rect -35 -318 -30 -312
rect -21 -318 -17 -312
rect 44 -317 49 -311
rect 58 -317 62 -311
rect 67 -317 72 -311
rect 81 -317 85 -311
rect 105 -317 110 -311
rect 119 -317 123 -311
rect 189 -316 194 -310
rect 203 -316 207 -310
rect 212 -316 217 -310
rect 226 -316 230 -310
rect 250 -316 255 -310
rect 264 -316 268 -310
rect 350 -319 355 -313
rect 364 -319 368 -313
rect 373 -319 378 -313
rect 387 -319 391 -313
rect 396 -319 401 -313
rect 410 -319 414 -313
rect 419 -319 424 -313
rect 433 -319 437 -313
<< polysilicon >>
rect -6 -142 44 -139
rect -6 -237 -3 -142
rect 18 -161 21 -157
rect 41 -161 44 -142
rect 149 -141 199 -138
rect 72 -161 75 -157
rect 95 -161 98 -157
rect 18 -206 21 -167
rect 41 -173 44 -167
rect 72 -185 75 -167
rect 95 -185 98 -167
rect 70 -189 75 -185
rect 88 -189 98 -185
rect 18 -209 44 -206
rect 18 -216 21 -212
rect 41 -216 44 -209
rect 72 -216 75 -189
rect 95 -216 98 -189
rect 18 -237 21 -220
rect 41 -224 44 -220
rect 72 -223 75 -220
rect 95 -222 98 -220
rect 83 -223 98 -222
rect 83 -224 94 -223
rect 41 -226 63 -224
rect 61 -228 63 -226
rect 83 -228 85 -224
rect 61 -230 85 -228
rect 114 -237 119 -189
rect -6 -240 119 -237
rect 149 -236 152 -141
rect 173 -160 176 -156
rect 196 -160 199 -141
rect 227 -160 230 -156
rect 250 -160 253 -156
rect 173 -205 176 -166
rect 196 -172 199 -166
rect 227 -184 230 -166
rect 250 -184 253 -166
rect 225 -188 230 -184
rect 243 -188 253 -184
rect 173 -208 199 -205
rect 173 -215 176 -211
rect 196 -215 199 -208
rect 227 -215 230 -188
rect 250 -215 253 -188
rect 173 -236 176 -219
rect 196 -223 199 -219
rect 227 -222 230 -219
rect 250 -221 253 -219
rect 238 -222 253 -221
rect 238 -223 249 -222
rect 196 -225 218 -223
rect 216 -227 218 -225
rect 238 -227 240 -223
rect 216 -229 240 -227
rect 269 -236 274 -188
rect 149 -239 274 -236
rect -88 -312 -85 -309
rect -65 -312 -62 -309
rect -27 -312 -24 -309
rect 52 -311 55 -308
rect 75 -311 78 -308
rect 113 -311 116 -308
rect 197 -310 200 -307
rect 220 -310 223 -307
rect 258 -310 261 -307
rect 358 -313 361 -309
rect 381 -313 384 -309
rect 404 -313 407 -309
rect 427 -313 430 -309
rect -88 -329 -85 -318
rect -90 -333 -85 -329
rect -88 -349 -85 -333
rect -65 -338 -62 -318
rect -27 -328 -24 -318
rect 52 -328 55 -317
rect -29 -332 -24 -328
rect 50 -332 55 -328
rect -67 -342 -62 -338
rect -65 -349 -62 -342
rect -27 -349 -24 -332
rect 52 -348 55 -332
rect 75 -337 78 -317
rect 113 -327 116 -317
rect 197 -327 200 -316
rect 111 -331 116 -327
rect 195 -331 200 -327
rect 73 -341 78 -337
rect 75 -348 78 -341
rect 113 -348 116 -331
rect 197 -347 200 -331
rect 220 -336 223 -316
rect 258 -326 261 -316
rect 256 -330 261 -326
rect 218 -340 223 -336
rect 220 -347 223 -340
rect 258 -347 261 -330
rect 358 -342 361 -319
rect 381 -342 384 -319
rect 404 -342 407 -319
rect 427 -331 430 -319
rect 425 -335 430 -331
rect 427 -342 430 -335
rect 358 -351 361 -347
rect -88 -358 -85 -354
rect -65 -358 -62 -354
rect -27 -358 -24 -354
rect 52 -357 55 -353
rect 75 -357 78 -353
rect 113 -357 116 -353
rect 197 -356 200 -352
rect 220 -356 223 -352
rect 258 -356 261 -352
rect 381 -363 384 -347
rect 404 -372 407 -347
rect 427 -351 430 -347
<< polycontact >>
rect 65 -189 70 -185
rect 114 -189 119 -185
rect 94 -227 99 -223
rect 220 -188 225 -184
rect 269 -188 274 -184
rect 249 -226 254 -222
rect -95 -333 -90 -329
rect -34 -332 -29 -328
rect 45 -332 50 -328
rect -72 -342 -67 -338
rect 106 -331 111 -327
rect 190 -331 195 -327
rect 68 -341 73 -337
rect 251 -330 256 -326
rect 353 -330 358 -326
rect 213 -340 218 -336
rect 420 -335 425 -331
rect 381 -367 386 -363
rect 403 -376 408 -372
<< metal1 >>
rect -208 -127 233 -122
rect -208 -290 -203 -127
rect 10 -136 59 -132
rect 10 -161 15 -136
rect -184 -257 -38 -253
rect -184 -363 -178 -257
rect -23 -270 -20 -190
rect 10 -216 15 -167
rect 24 -151 46 -146
rect 24 -161 28 -151
rect 47 -161 51 -151
rect 24 -216 28 -167
rect 33 -216 38 -167
rect 47 -216 51 -167
rect 56 -185 59 -136
rect 71 -144 74 -127
rect 170 -135 214 -131
rect 64 -149 92 -144
rect 64 -161 69 -149
rect 87 -161 92 -149
rect 165 -160 170 -136
rect 59 -189 65 -185
rect 78 -194 82 -167
rect 56 -198 82 -194
rect 33 -228 38 -220
rect 56 -228 59 -198
rect 78 -216 82 -198
rect 101 -185 105 -167
rect 101 -189 114 -185
rect 101 -216 105 -189
rect 33 -231 59 -228
rect 165 -215 170 -166
rect 179 -150 206 -145
rect 179 -160 183 -150
rect 202 -160 206 -150
rect 179 -215 183 -166
rect 188 -215 193 -166
rect 202 -215 206 -166
rect 211 -184 214 -135
rect 230 -143 233 -127
rect 219 -148 247 -143
rect 219 -160 224 -148
rect 242 -160 247 -148
rect 211 -188 220 -184
rect 233 -193 237 -166
rect 211 -197 237 -193
rect 64 -231 68 -220
rect 87 -231 91 -220
rect 188 -227 193 -219
rect 211 -227 214 -197
rect 233 -215 237 -197
rect 256 -184 260 -166
rect 256 -188 269 -184
rect 256 -215 260 -188
rect 64 -235 91 -231
rect 76 -253 79 -235
rect 95 -241 98 -227
rect 188 -230 214 -227
rect 219 -230 223 -219
rect 242 -230 246 -219
rect 219 -234 246 -230
rect 233 -253 236 -234
rect 9 -257 236 -253
rect 250 -262 253 -226
rect 29 -266 253 -262
rect -136 -274 148 -270
rect -136 -329 -130 -274
rect -119 -281 -114 -280
rect -119 -284 94 -281
rect -119 -285 -114 -284
rect -118 -317 -115 -285
rect -71 -302 -68 -295
rect -103 -306 -9 -302
rect -96 -312 -91 -306
rect -73 -312 -68 -306
rect -35 -312 -30 -306
rect -82 -328 -78 -318
rect -59 -328 -55 -318
rect -21 -328 -17 -318
rect -136 -333 -95 -329
rect -82 -332 -34 -328
rect -21 -332 -8 -328
rect -114 -342 -72 -338
rect -59 -349 -55 -332
rect -21 -349 -17 -332
rect -78 -354 -73 -349
rect -96 -363 -92 -354
rect -35 -363 -31 -354
rect -184 -366 -35 -363
rect -184 -368 -178 -366
rect -11 -384 -8 -332
rect 2 -337 7 -284
rect 25 -328 28 -292
rect 60 -301 63 -295
rect 37 -305 131 -301
rect 44 -311 49 -305
rect 67 -311 72 -305
rect 105 -311 110 -305
rect 58 -327 62 -317
rect 81 -327 85 -317
rect 119 -327 123 -317
rect 25 -332 45 -328
rect 58 -331 106 -327
rect 119 -331 130 -327
rect 2 -341 68 -337
rect 81 -348 85 -331
rect 119 -348 123 -331
rect 62 -353 67 -348
rect 44 -362 48 -353
rect 105 -361 109 -353
rect 44 -363 105 -362
rect 48 -365 105 -363
rect 127 -372 130 -331
rect 141 -336 148 -274
rect 163 -327 169 -266
rect 206 -294 369 -291
rect 202 -300 205 -295
rect 182 -304 276 -300
rect 364 -301 369 -294
rect 189 -310 194 -304
rect 212 -310 217 -304
rect 250 -310 255 -304
rect 350 -305 424 -301
rect 203 -326 207 -316
rect 226 -326 230 -316
rect 264 -326 268 -316
rect 350 -313 355 -305
rect 419 -313 424 -305
rect 368 -319 373 -313
rect 391 -319 396 -313
rect 163 -331 190 -327
rect 203 -330 251 -326
rect 264 -330 353 -326
rect 141 -340 213 -336
rect 226 -347 230 -330
rect 264 -347 268 -330
rect 410 -331 414 -319
rect 433 -331 437 -319
rect 410 -335 420 -331
rect 433 -335 442 -331
rect 410 -336 414 -335
rect 364 -339 414 -336
rect 364 -342 368 -339
rect 387 -342 391 -339
rect 410 -342 414 -339
rect 433 -342 437 -335
rect 207 -352 212 -347
rect 189 -360 193 -352
rect 250 -360 254 -352
rect 350 -354 354 -347
rect 373 -354 377 -347
rect 396 -354 400 -347
rect 419 -354 423 -347
rect 350 -355 423 -354
rect 270 -358 423 -355
rect 270 -360 275 -358
rect 250 -361 275 -360
rect 193 -364 275 -361
rect 279 -367 381 -364
rect 279 -372 283 -367
rect 127 -376 283 -372
rect 292 -376 403 -372
rect 292 -384 295 -376
rect -11 -389 295 -384
<< m2contact >>
rect -24 -190 -19 -185
rect -208 -295 -203 -290
rect -38 -257 -33 -252
rect 46 -151 51 -146
rect 165 -136 170 -131
rect 54 -190 59 -185
rect 4 -257 9 -252
rect 94 -246 99 -241
rect 24 -266 29 -261
rect 94 -284 99 -279
rect -72 -295 -67 -290
rect -119 -322 -114 -317
rect -119 -343 -114 -338
rect -35 -368 -30 -363
rect 24 -292 29 -287
rect 59 -295 64 -290
rect 43 -368 48 -363
rect 105 -366 110 -361
rect 201 -295 206 -290
rect 188 -365 193 -360
<< metal2 >>
rect 126 -135 165 -131
rect 126 -138 129 -135
rect 47 -142 129 -138
rect 47 -146 50 -142
rect -19 -189 54 -186
rect -33 -256 4 -253
rect 25 -287 28 -266
rect 95 -279 98 -246
rect -203 -294 -72 -291
rect -67 -294 14 -291
rect 11 -297 14 -294
rect 38 -294 59 -291
rect 38 -297 41 -294
rect 64 -294 201 -291
rect 11 -300 41 -297
rect -118 -338 -115 -322
rect -30 -367 43 -364
rect 110 -365 188 -362
<< labels >>
rlabel metal1 148 -126 153 -123 5 vdd
rlabel polysilicon 245 -187 249 -185 1 C
rlabel polysilicon 71 -188 75 -186 1 A
rlabel polysilicon 91 -188 95 -186 1 B
rlabel metal1 189 -149 193 -147 1 sum
rlabel metal1 161 -257 166 -255 1 gnd
rlabel metal1 438 -334 441 -332 7 carry
<< end >>
