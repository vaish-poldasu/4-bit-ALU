magic
tech scmos
timestamp 1700213876
<< nwell >>
rect 44 32 98 50
rect 110 32 141 50
rect 152 32 206 50
rect 218 32 249 50
rect 264 32 318 50
rect 330 32 361 50
rect 376 32 430 50
rect 442 32 473 50
rect 487 32 541 50
rect 553 32 584 50
rect 599 32 653 50
rect 665 32 696 50
rect 711 32 765 50
rect 777 32 808 50
rect 823 32 877 50
rect 889 32 920 50
<< ntransistor >>
rect 59 2 62 7
rect 82 2 85 7
rect 125 2 128 7
rect 167 2 170 7
rect 190 2 193 7
rect 233 2 236 7
rect 279 2 282 7
rect 302 2 305 7
rect 345 2 348 7
rect 391 2 394 7
rect 414 2 417 7
rect 457 2 460 7
rect 502 2 505 7
rect 525 2 528 7
rect 568 2 571 7
rect 614 2 617 7
rect 637 2 640 7
rect 680 2 683 7
rect 726 2 729 7
rect 749 2 752 7
rect 792 2 795 7
rect 838 2 841 7
rect 861 2 864 7
rect 904 2 907 7
<< ptransistor >>
rect 59 38 62 44
rect 82 38 85 44
rect 125 38 128 44
rect 167 38 170 44
rect 190 38 193 44
rect 233 38 236 44
rect 279 38 282 44
rect 302 38 305 44
rect 345 38 348 44
rect 391 38 394 44
rect 414 38 417 44
rect 457 38 460 44
rect 502 38 505 44
rect 525 38 528 44
rect 568 38 571 44
rect 614 38 617 44
rect 637 38 640 44
rect 680 38 683 44
rect 726 38 729 44
rect 749 38 752 44
rect 792 38 795 44
rect 838 38 841 44
rect 861 38 864 44
rect 904 38 907 44
<< ndiffusion >>
rect 55 2 59 7
rect 62 2 65 7
rect 78 2 82 7
rect 85 2 88 7
rect 121 2 125 7
rect 128 2 131 7
rect 163 2 167 7
rect 170 2 173 7
rect 186 2 190 7
rect 193 2 196 7
rect 229 2 233 7
rect 236 2 239 7
rect 275 2 279 7
rect 282 2 285 7
rect 298 2 302 7
rect 305 2 308 7
rect 341 2 345 7
rect 348 2 351 7
rect 387 2 391 7
rect 394 2 397 7
rect 410 2 414 7
rect 417 2 420 7
rect 453 2 457 7
rect 460 2 463 7
rect 498 2 502 7
rect 505 2 508 7
rect 521 2 525 7
rect 528 2 531 7
rect 564 2 568 7
rect 571 2 574 7
rect 610 2 614 7
rect 617 2 620 7
rect 633 2 637 7
rect 640 2 643 7
rect 676 2 680 7
rect 683 2 686 7
rect 722 2 726 7
rect 729 2 732 7
rect 745 2 749 7
rect 752 2 755 7
rect 788 2 792 7
rect 795 2 798 7
rect 834 2 838 7
rect 841 2 844 7
rect 857 2 861 7
rect 864 2 867 7
rect 900 2 904 7
rect 907 2 910 7
<< pdiffusion >>
rect 56 38 59 44
rect 62 38 65 44
rect 79 38 82 44
rect 85 38 88 44
rect 122 38 125 44
rect 128 38 131 44
rect 164 38 167 44
rect 170 38 173 44
rect 187 38 190 44
rect 193 38 196 44
rect 230 38 233 44
rect 236 38 239 44
rect 276 38 279 44
rect 282 38 285 44
rect 299 38 302 44
rect 305 38 308 44
rect 342 38 345 44
rect 348 38 351 44
rect 388 38 391 44
rect 394 38 397 44
rect 411 38 414 44
rect 417 38 420 44
rect 454 38 457 44
rect 460 38 463 44
rect 499 38 502 44
rect 505 38 508 44
rect 522 38 525 44
rect 528 38 531 44
rect 565 38 568 44
rect 571 38 574 44
rect 611 38 614 44
rect 617 38 620 44
rect 634 38 637 44
rect 640 38 643 44
rect 677 38 680 44
rect 683 38 686 44
rect 723 38 726 44
rect 729 38 732 44
rect 746 38 749 44
rect 752 38 755 44
rect 789 38 792 44
rect 795 38 798 44
rect 835 38 838 44
rect 841 38 844 44
rect 858 38 861 44
rect 864 38 867 44
rect 901 38 904 44
rect 907 38 910 44
<< ndcontact >>
rect 51 2 55 7
rect 65 2 69 7
rect 74 2 78 7
rect 88 2 92 7
rect 117 2 121 7
rect 131 2 135 7
rect 159 2 163 7
rect 173 2 177 7
rect 182 2 186 7
rect 196 2 200 7
rect 225 2 229 7
rect 239 2 243 7
rect 271 2 275 7
rect 285 2 289 7
rect 294 2 298 7
rect 308 2 312 7
rect 337 2 341 7
rect 351 2 355 7
rect 383 2 387 7
rect 397 2 401 7
rect 406 2 410 7
rect 420 2 424 7
rect 449 2 453 7
rect 463 2 467 7
rect 494 2 498 7
rect 508 2 512 7
rect 517 2 521 7
rect 531 2 535 7
rect 560 2 564 7
rect 574 2 578 7
rect 606 2 610 7
rect 620 2 624 7
rect 629 2 633 7
rect 643 2 647 7
rect 672 2 676 7
rect 686 2 690 7
rect 718 2 722 7
rect 732 2 736 7
rect 741 2 745 7
rect 755 2 759 7
rect 784 2 788 7
rect 798 2 802 7
rect 830 2 834 7
rect 844 2 848 7
rect 853 2 857 7
rect 867 2 871 7
rect 896 2 900 7
rect 910 2 914 7
<< pdcontact >>
rect 51 38 56 44
rect 65 38 69 44
rect 74 38 79 44
rect 88 38 92 44
rect 117 38 122 44
rect 131 38 135 44
rect 159 38 164 44
rect 173 38 177 44
rect 182 38 187 44
rect 196 38 200 44
rect 225 38 230 44
rect 239 38 243 44
rect 271 38 276 44
rect 285 38 289 44
rect 294 38 299 44
rect 308 38 312 44
rect 337 38 342 44
rect 351 38 355 44
rect 383 38 388 44
rect 397 38 401 44
rect 406 38 411 44
rect 420 38 424 44
rect 449 38 454 44
rect 463 38 467 44
rect 494 38 499 44
rect 508 38 512 44
rect 517 38 522 44
rect 531 38 535 44
rect 560 38 565 44
rect 574 38 578 44
rect 606 38 611 44
rect 620 38 624 44
rect 629 38 634 44
rect 643 38 647 44
rect 672 38 677 44
rect 686 38 690 44
rect 718 38 723 44
rect 732 38 736 44
rect 741 38 746 44
rect 755 38 759 44
rect 784 38 789 44
rect 798 38 802 44
rect 830 38 835 44
rect 844 38 848 44
rect 853 38 858 44
rect 867 38 871 44
rect 896 38 901 44
rect 910 38 914 44
<< polysilicon >>
rect 59 44 62 63
rect 82 44 85 47
rect 125 44 128 47
rect 167 44 170 63
rect 190 44 193 47
rect 233 44 236 47
rect 279 44 282 63
rect 302 44 305 47
rect 345 44 348 47
rect 391 44 394 63
rect 414 44 417 47
rect 457 44 460 47
rect 502 44 505 63
rect 525 44 528 47
rect 568 44 571 47
rect 614 44 617 63
rect 637 44 640 47
rect 680 44 683 47
rect 726 44 729 63
rect 749 44 752 47
rect 792 44 795 47
rect 838 44 841 63
rect 861 44 864 47
rect 904 44 907 47
rect 59 7 62 38
rect 82 7 85 38
rect 125 28 128 38
rect 123 24 128 28
rect 125 7 128 24
rect 167 7 170 38
rect 190 7 193 38
rect 233 28 236 38
rect 231 24 236 28
rect 233 7 236 24
rect 279 7 282 38
rect 302 7 305 38
rect 345 28 348 38
rect 343 24 348 28
rect 345 7 348 24
rect 391 7 394 38
rect 414 7 417 38
rect 457 28 460 38
rect 455 24 460 28
rect 457 7 460 24
rect 502 7 505 38
rect 525 7 528 38
rect 568 28 571 38
rect 566 24 571 28
rect 568 7 571 24
rect 614 7 617 38
rect 637 7 640 38
rect 680 28 683 38
rect 678 24 683 28
rect 680 7 683 24
rect 726 7 729 38
rect 749 7 752 38
rect 792 28 795 38
rect 790 24 795 28
rect 792 7 795 24
rect 838 7 841 38
rect 861 7 864 38
rect 904 28 907 38
rect 902 24 907 28
rect 904 7 907 24
rect 59 -2 62 2
rect 82 -2 85 2
rect 125 -2 128 2
rect 167 -2 170 2
rect 190 -2 193 2
rect 233 -2 236 2
rect 279 -2 282 2
rect 302 -2 305 2
rect 345 -2 348 2
rect 391 -2 394 2
rect 414 -2 417 2
rect 457 -2 460 2
rect 502 -2 505 2
rect 525 -2 528 2
rect 568 -2 571 2
rect 614 -2 617 2
rect 637 -2 640 2
rect 680 -2 683 2
rect 726 -2 729 2
rect 749 -2 752 2
rect 792 -2 795 2
rect 838 -2 841 2
rect 861 -2 864 2
rect 904 -2 907 2
<< polycontact >>
rect 58 63 63 67
rect 166 63 171 67
rect 278 63 283 67
rect 390 63 395 67
rect 501 63 506 67
rect 613 63 618 67
rect 725 63 730 67
rect 837 63 842 67
rect 118 24 123 28
rect 226 24 231 28
rect 338 24 343 28
rect 450 24 455 28
rect 561 24 566 28
rect 673 24 678 28
rect 785 24 790 28
rect 897 24 902 28
<< metal1 >>
rect 58 67 63 83
rect 63 63 166 66
rect 171 63 278 66
rect 283 63 390 66
rect 395 63 501 66
rect 506 63 613 66
rect 618 63 725 66
rect 730 63 837 66
rect 44 50 920 54
rect 51 44 56 50
rect 74 44 79 50
rect 117 44 122 50
rect 159 44 164 50
rect 182 44 187 50
rect 225 44 230 50
rect 271 44 276 50
rect 294 44 299 50
rect 337 44 342 50
rect 383 44 388 50
rect 406 44 411 50
rect 449 44 454 50
rect 494 44 499 50
rect 517 44 522 50
rect 560 44 565 50
rect 606 44 611 50
rect 629 44 634 50
rect 672 44 677 50
rect 718 44 723 50
rect 741 44 746 50
rect 784 44 789 50
rect 830 44 835 50
rect 853 44 858 50
rect 896 44 901 50
rect 65 28 69 38
rect 88 28 92 38
rect 131 28 135 38
rect 173 28 177 38
rect 196 28 200 38
rect 239 28 243 38
rect 285 28 289 38
rect 308 28 312 38
rect 351 28 355 38
rect 397 28 401 38
rect 420 28 424 38
rect 463 28 467 38
rect 508 28 512 38
rect 531 28 535 38
rect 574 28 578 38
rect 620 28 624 38
rect 643 28 647 38
rect 686 28 690 38
rect 732 28 736 38
rect 755 28 759 38
rect 798 28 802 38
rect 844 28 848 38
rect 867 28 871 38
rect 910 28 914 38
rect 65 24 118 28
rect 131 24 141 28
rect 173 24 226 28
rect 239 24 249 28
rect 285 24 338 28
rect 351 24 361 28
rect 397 24 450 28
rect 463 24 473 28
rect 508 24 561 28
rect 574 24 584 28
rect 620 24 673 28
rect 686 24 696 28
rect 732 24 785 28
rect 798 24 808 28
rect 844 24 897 28
rect 910 24 920 28
rect 88 7 92 24
rect 131 7 135 24
rect 196 7 200 24
rect 239 7 243 24
rect 308 7 312 24
rect 351 7 355 24
rect 420 7 424 24
rect 463 7 467 24
rect 531 7 535 24
rect 574 7 578 24
rect 643 7 647 24
rect 686 7 690 24
rect 755 7 759 24
rect 798 7 802 24
rect 867 7 871 24
rect 910 7 914 24
rect 69 2 74 7
rect 177 2 182 7
rect 289 2 294 7
rect 401 2 406 7
rect 512 2 517 7
rect 624 2 629 7
rect 736 2 741 7
rect 848 2 853 7
rect 51 -7 55 2
rect 117 -6 121 2
rect 159 -6 163 2
rect 117 -7 163 -6
rect 225 -6 229 2
rect 271 -6 275 2
rect 225 -7 275 -6
rect 337 -6 341 2
rect 383 -6 387 2
rect 337 -7 387 -6
rect 449 -6 453 2
rect 494 -6 498 2
rect 449 -7 498 -6
rect 560 -6 564 2
rect 606 -6 610 2
rect 560 -7 610 -6
rect 672 -6 676 2
rect 718 -6 722 2
rect 672 -7 722 -6
rect 784 -6 788 2
rect 830 -6 834 2
rect 784 -7 834 -6
rect 896 -7 900 2
rect 51 -10 900 -7
<< labels >>
rlabel metal1 62 -10 65 -8 1 gnd
rlabel metal1 68 51 71 53 5 vdd
rlabel metal1 58 70 62 73 1 en
rlabel polysilicon 82 18 85 21 1 B3
rlabel polysilicon 190 19 193 22 1 B2
rlabel polysilicon 302 19 305 22 1 B1
rlabel polysilicon 414 19 417 22 1 B0
rlabel polysilicon 525 20 528 23 1 A3
rlabel polysilicon 637 19 640 22 1 A2
rlabel polysilicon 749 20 752 23 1 A1
rlabel polysilicon 861 20 864 23 1 A0
rlabel metal1 915 25 918 28 7 A0_out
rlabel metal1 802 25 805 28 1 A1_out
rlabel metal1 691 24 694 27 1 A2_out
rlabel metal1 578 24 581 27 1 A3_out
rlabel metal1 468 24 471 27 1 B0_out
rlabel metal1 356 24 359 27 1 B1_out
rlabel metal1 244 24 247 27 1 B2_out
rlabel metal1 136 24 139 27 1 B3_out
<< end >>
