magic
tech scmos
timestamp 1699895379
<< nwell >>
rect 174 157 228 175
rect 235 157 266 175
rect 322 174 353 192
rect 412 161 466 179
rect 473 161 504 179
rect 543 161 597 179
rect 604 161 635 179
rect 699 161 753 179
rect 760 161 791 179
rect 321 106 352 124
<< ntransistor >>
rect 337 154 340 159
rect 189 127 192 132
rect 212 127 215 132
rect 250 127 253 132
rect 427 131 430 136
rect 450 131 453 136
rect 488 131 491 136
rect 558 131 561 136
rect 581 131 584 136
rect 619 131 622 136
rect 714 131 717 136
rect 737 131 740 136
rect 775 131 778 136
rect 336 86 339 91
<< ptransistor >>
rect 337 180 340 186
rect 189 163 192 169
rect 212 163 215 169
rect 250 163 253 169
rect 427 167 430 173
rect 450 167 453 173
rect 488 167 491 173
rect 558 167 561 173
rect 581 167 584 173
rect 619 167 622 173
rect 714 167 717 173
rect 737 167 740 173
rect 775 167 778 173
rect 336 112 339 118
<< ndiffusion >>
rect 333 154 337 159
rect 340 154 343 159
rect 185 127 189 132
rect 192 127 195 132
rect 208 127 212 132
rect 215 127 218 132
rect 246 127 250 132
rect 253 127 256 132
rect 423 131 427 136
rect 430 131 433 136
rect 446 131 450 136
rect 453 131 456 136
rect 484 131 488 136
rect 491 131 494 136
rect 554 131 558 136
rect 561 131 564 136
rect 577 131 581 136
rect 584 131 587 136
rect 615 131 619 136
rect 622 131 625 136
rect 710 131 714 136
rect 717 131 720 136
rect 733 131 737 136
rect 740 131 743 136
rect 771 131 775 136
rect 778 131 781 136
rect 332 86 336 91
rect 339 86 342 91
<< pdiffusion >>
rect 334 180 337 186
rect 340 180 343 186
rect 186 163 189 169
rect 192 163 195 169
rect 209 163 212 169
rect 215 163 218 169
rect 247 163 250 169
rect 253 163 256 169
rect 424 167 427 173
rect 430 167 433 173
rect 447 167 450 173
rect 453 167 456 173
rect 485 167 488 173
rect 491 167 494 173
rect 555 167 558 173
rect 561 167 564 173
rect 578 167 581 173
rect 584 167 587 173
rect 616 167 619 173
rect 622 167 625 173
rect 711 167 714 173
rect 717 167 720 173
rect 734 167 737 173
rect 740 167 743 173
rect 772 167 775 173
rect 778 167 781 173
rect 333 112 336 118
rect 339 112 342 118
<< ndcontact >>
rect 329 154 333 159
rect 343 154 347 159
rect 181 127 185 132
rect 195 127 199 132
rect 204 127 208 132
rect 218 127 222 132
rect 242 127 246 132
rect 256 127 260 132
rect 419 131 423 136
rect 433 131 437 136
rect 442 131 446 136
rect 456 131 460 136
rect 480 131 484 136
rect 494 131 498 136
rect 550 131 554 136
rect 564 131 568 136
rect 573 131 577 136
rect 587 131 591 136
rect 611 131 615 136
rect 625 131 629 136
rect 706 131 710 136
rect 720 131 724 136
rect 729 131 733 136
rect 743 131 747 136
rect 767 131 771 136
rect 781 131 785 136
rect 328 86 332 91
rect 342 86 346 91
<< pdcontact >>
rect 329 180 334 186
rect 343 180 347 186
rect 181 163 186 169
rect 195 163 199 169
rect 204 163 209 169
rect 218 163 222 169
rect 242 163 247 169
rect 256 163 260 169
rect 419 167 424 173
rect 433 167 437 173
rect 442 167 447 173
rect 456 167 460 173
rect 480 167 485 173
rect 494 167 498 173
rect 550 167 555 173
rect 564 167 568 173
rect 573 167 578 173
rect 587 167 591 173
rect 611 167 616 173
rect 625 167 629 173
rect 706 167 711 173
rect 720 167 724 173
rect 729 167 734 173
rect 743 167 747 173
rect 767 167 772 173
rect 781 167 785 173
rect 328 112 333 118
rect 342 112 346 118
<< polysilicon >>
rect 337 186 340 189
rect 189 169 192 172
rect 212 169 215 172
rect 250 169 253 172
rect 337 169 340 180
rect 427 173 430 176
rect 450 173 453 176
rect 488 173 491 176
rect 558 173 561 176
rect 581 173 584 176
rect 619 173 622 176
rect 714 173 717 176
rect 737 173 740 176
rect 775 173 778 176
rect 335 165 340 169
rect 189 132 192 163
rect 212 142 215 163
rect 250 153 253 163
rect 337 159 340 165
rect 427 156 430 167
rect 248 149 253 153
rect 210 138 215 142
rect 212 132 215 138
rect 250 132 253 149
rect 337 147 340 154
rect 425 152 430 156
rect 427 136 430 152
rect 450 147 453 167
rect 488 157 491 167
rect 486 153 491 157
rect 558 156 561 167
rect 448 143 453 147
rect 450 136 453 143
rect 488 136 491 153
rect 556 152 561 156
rect 558 136 561 152
rect 581 147 584 167
rect 619 157 622 167
rect 617 153 622 157
rect 714 156 717 167
rect 579 143 584 147
rect 581 136 584 143
rect 619 136 622 153
rect 712 152 717 156
rect 714 136 717 152
rect 737 147 740 167
rect 775 157 778 167
rect 773 153 778 157
rect 735 143 740 147
rect 737 136 740 143
rect 775 136 778 153
rect 427 127 430 131
rect 450 127 453 131
rect 488 127 491 131
rect 558 127 561 131
rect 581 127 584 131
rect 619 127 622 131
rect 714 127 717 131
rect 737 127 740 131
rect 775 127 778 131
rect 189 123 192 127
rect 212 123 215 127
rect 250 123 253 127
rect 336 118 339 121
rect 336 101 339 112
rect 334 97 339 101
rect 336 91 339 97
rect 336 79 339 86
<< polycontact >>
rect 330 165 335 169
rect 184 147 189 151
rect 243 149 248 153
rect 205 138 210 142
rect 420 152 425 156
rect 481 153 486 157
rect 443 143 448 147
rect 551 152 556 156
rect 612 153 617 157
rect 574 143 579 147
rect 707 152 712 156
rect 768 153 773 157
rect 730 143 735 147
rect 329 97 334 101
<< metal1 >>
rect 312 220 680 223
rect 161 187 291 190
rect 161 151 164 187
rect 174 175 261 179
rect 181 169 186 175
rect 204 169 209 175
rect 242 169 247 175
rect 288 169 291 187
rect 312 169 315 220
rect 364 201 528 204
rect 327 192 353 197
rect 329 186 334 192
rect 343 169 347 180
rect 364 169 367 201
rect 454 183 459 191
rect 412 179 504 183
rect 288 165 330 169
rect 343 165 367 169
rect 419 173 424 179
rect 442 173 447 179
rect 480 173 485 179
rect 195 153 199 163
rect 218 153 222 163
rect 256 153 260 163
rect 343 159 347 165
rect 364 156 367 165
rect 433 157 437 167
rect 456 157 460 167
rect 494 157 498 167
rect 161 147 184 151
rect 195 149 243 153
rect 256 149 266 153
rect 161 138 205 142
rect 161 101 164 138
rect 218 132 222 149
rect 256 132 260 149
rect 329 146 333 154
rect 364 152 420 156
rect 433 153 481 157
rect 494 153 504 157
rect 524 156 528 201
rect 590 183 595 191
rect 543 179 635 183
rect 550 173 555 179
rect 573 173 578 179
rect 611 173 616 179
rect 564 157 568 167
rect 587 157 591 167
rect 625 157 629 167
rect 321 143 353 146
rect 364 143 443 147
rect 199 127 204 132
rect 181 118 185 127
rect 242 118 246 127
rect 321 124 352 129
rect 181 115 246 118
rect 328 118 333 124
rect 342 101 346 112
rect 364 101 367 143
rect 456 136 460 153
rect 494 136 498 153
rect 524 152 551 156
rect 564 153 612 157
rect 625 153 635 157
rect 677 156 680 220
rect 728 183 733 191
rect 699 179 791 183
rect 706 173 711 179
rect 729 173 734 179
rect 767 173 772 179
rect 720 157 724 167
rect 743 157 747 167
rect 781 157 785 167
rect 548 143 574 147
rect 587 136 591 153
rect 625 136 629 153
rect 677 152 707 156
rect 720 153 768 157
rect 781 153 791 157
rect 437 131 442 136
rect 568 131 573 136
rect 678 143 730 147
rect 419 122 423 131
rect 480 122 484 131
rect 419 119 484 122
rect 550 122 554 131
rect 611 122 615 131
rect 550 119 615 122
rect 161 97 329 101
rect 342 97 367 101
rect 447 102 451 119
rect 577 102 581 119
rect 379 99 664 102
rect 306 70 309 97
rect 342 91 346 97
rect 364 87 367 97
rect 678 87 681 143
rect 743 136 747 153
rect 781 136 785 153
rect 724 131 729 136
rect 706 122 710 131
rect 767 122 771 131
rect 706 119 771 122
rect 742 102 746 119
rect 696 99 746 102
rect 328 78 332 86
rect 364 84 681 87
rect 321 75 351 78
rect 306 67 523 70
<< m2contact >>
rect 261 175 266 180
rect 322 192 327 197
rect 353 192 358 197
rect 454 191 459 196
rect 316 143 321 148
rect 590 191 595 196
rect 352 124 357 129
rect 246 114 251 119
rect 728 191 733 196
rect 543 142 548 147
rect 374 98 379 103
rect 664 98 669 103
rect 691 98 696 103
rect 316 75 321 80
rect 351 75 356 80
rect 523 67 528 72
<< metal2 >>
rect 263 193 322 196
rect 263 180 266 193
rect 358 193 454 196
rect 316 118 319 143
rect 354 129 357 192
rect 459 193 590 196
rect 595 193 728 196
rect 733 193 734 196
rect 523 143 543 147
rect 251 115 319 118
rect 316 80 319 115
rect 374 78 377 98
rect 356 75 377 78
rect 523 72 526 143
rect 669 99 691 102
<< labels >>
rlabel metal1 338 193 341 195 1 vdd
rlabel metal1 335 75 339 77 1 gnd
rlabel metal1 260 150 264 152 1 D3
rlabel metal1 786 154 790 156 7 D2
rlabel metal1 630 154 634 156 1 D1
rlabel metal1 498 154 502 156 1 D0
rlabel metal1 321 98 325 100 1 S0
rlabel metal1 322 166 326 168 1 S1
<< end >>
