magic
tech scmos
timestamp 1700211523
<< nwell >>
rect -480 -842 -372 -824
rect 310 -842 418 -824
rect 1292 -842 1400 -824
rect 2176 -842 2284 -824
rect -467 -1153 -359 -1135
rect -312 -1152 -204 -1134
rect 334 -1151 442 -1133
rect 489 -1150 597 -1132
rect 1237 -1151 1345 -1133
rect 1392 -1150 1500 -1132
rect 2105 -1150 2213 -1132
rect 2260 -1149 2368 -1131
rect -573 -1304 -519 -1286
rect -512 -1304 -481 -1286
rect -433 -1303 -379 -1285
rect -372 -1303 -341 -1285
rect -288 -1302 -234 -1284
rect -227 -1302 -196 -1284
rect -127 -1305 -27 -1287
rect 228 -1302 282 -1284
rect 289 -1302 320 -1284
rect 368 -1301 422 -1283
rect 429 -1301 460 -1283
rect 513 -1300 567 -1282
rect 574 -1300 605 -1282
rect 674 -1303 774 -1285
rect 1131 -1302 1185 -1284
rect 1192 -1302 1223 -1284
rect 1271 -1301 1325 -1283
rect 1332 -1301 1363 -1283
rect 1416 -1300 1470 -1282
rect 1477 -1300 1508 -1282
rect 1577 -1303 1677 -1285
rect 1999 -1301 2053 -1283
rect 2060 -1301 2091 -1283
rect 2139 -1300 2193 -1282
rect 2200 -1300 2231 -1282
rect 2284 -1299 2338 -1281
rect 2345 -1299 2376 -1281
rect 2445 -1302 2545 -1284
<< ntransistor >>
rect -465 -889 -462 -885
rect -442 -889 -439 -885
rect -411 -889 -408 -885
rect -388 -889 -385 -885
rect 325 -889 328 -885
rect 348 -889 351 -885
rect 379 -889 382 -885
rect 402 -889 405 -885
rect 1307 -889 1310 -885
rect 1330 -889 1333 -885
rect 1361 -889 1364 -885
rect 1384 -889 1387 -885
rect 2191 -889 2194 -885
rect 2214 -889 2217 -885
rect 2245 -889 2248 -885
rect 2268 -889 2271 -885
rect -452 -1200 -449 -1196
rect -429 -1200 -426 -1196
rect -398 -1200 -395 -1196
rect -375 -1200 -372 -1196
rect -297 -1199 -294 -1195
rect -274 -1199 -271 -1195
rect -243 -1199 -240 -1195
rect -220 -1199 -217 -1195
rect 349 -1198 352 -1194
rect 372 -1198 375 -1194
rect 403 -1198 406 -1194
rect 426 -1198 429 -1194
rect 504 -1197 507 -1193
rect 527 -1197 530 -1193
rect 558 -1197 561 -1193
rect 581 -1197 584 -1193
rect 1252 -1198 1255 -1194
rect 1275 -1198 1278 -1194
rect 1306 -1198 1309 -1194
rect 1329 -1198 1332 -1194
rect 1407 -1197 1410 -1193
rect 1430 -1197 1433 -1193
rect 1461 -1197 1464 -1193
rect 1484 -1197 1487 -1193
rect 2120 -1197 2123 -1193
rect 2143 -1197 2146 -1193
rect 2174 -1197 2177 -1193
rect 2197 -1197 2200 -1193
rect 2275 -1196 2278 -1192
rect 2298 -1196 2301 -1192
rect 2329 -1196 2332 -1192
rect 2352 -1196 2355 -1192
rect -112 -1327 -109 -1322
rect -89 -1327 -86 -1322
rect -66 -1327 -63 -1322
rect -43 -1327 -40 -1322
rect 689 -1325 692 -1320
rect 712 -1325 715 -1320
rect 735 -1325 738 -1320
rect 758 -1325 761 -1320
rect -558 -1334 -555 -1329
rect -535 -1334 -532 -1329
rect -497 -1334 -494 -1329
rect -418 -1333 -415 -1328
rect -395 -1333 -392 -1328
rect -357 -1333 -354 -1328
rect -273 -1332 -270 -1327
rect -250 -1332 -247 -1327
rect -212 -1332 -209 -1327
rect 243 -1332 246 -1327
rect 266 -1332 269 -1327
rect 304 -1332 307 -1327
rect 383 -1331 386 -1326
rect 406 -1331 409 -1326
rect 444 -1331 447 -1326
rect 528 -1330 531 -1325
rect 551 -1330 554 -1325
rect 589 -1330 592 -1325
rect 1592 -1325 1595 -1320
rect 1615 -1325 1618 -1320
rect 1638 -1325 1641 -1320
rect 1661 -1325 1664 -1320
rect 1146 -1332 1149 -1327
rect 1169 -1332 1172 -1327
rect 1207 -1332 1210 -1327
rect 1286 -1331 1289 -1326
rect 1309 -1331 1312 -1326
rect 1347 -1331 1350 -1326
rect 1431 -1330 1434 -1325
rect 1454 -1330 1457 -1325
rect 1492 -1330 1495 -1325
rect 2460 -1324 2463 -1319
rect 2483 -1324 2486 -1319
rect 2506 -1324 2509 -1319
rect 2529 -1324 2532 -1319
rect 2014 -1331 2017 -1326
rect 2037 -1331 2040 -1326
rect 2075 -1331 2078 -1326
rect 2154 -1330 2157 -1325
rect 2177 -1330 2180 -1325
rect 2215 -1330 2218 -1325
rect 2299 -1329 2302 -1324
rect 2322 -1329 2325 -1324
rect 2360 -1329 2363 -1324
<< ptransistor >>
rect -465 -836 -462 -830
rect -442 -836 -439 -830
rect -411 -836 -408 -830
rect -388 -836 -385 -830
rect 325 -836 328 -830
rect 348 -836 351 -830
rect 379 -836 382 -830
rect 402 -836 405 -830
rect 1307 -836 1310 -830
rect 1330 -836 1333 -830
rect 1361 -836 1364 -830
rect 1384 -836 1387 -830
rect 2191 -836 2194 -830
rect 2214 -836 2217 -830
rect 2245 -836 2248 -830
rect 2268 -836 2271 -830
rect -452 -1147 -449 -1141
rect -429 -1147 -426 -1141
rect -398 -1147 -395 -1141
rect -375 -1147 -372 -1141
rect -297 -1146 -294 -1140
rect -274 -1146 -271 -1140
rect -243 -1146 -240 -1140
rect -220 -1146 -217 -1140
rect 349 -1145 352 -1139
rect 372 -1145 375 -1139
rect 403 -1145 406 -1139
rect 426 -1145 429 -1139
rect 504 -1144 507 -1138
rect 527 -1144 530 -1138
rect 558 -1144 561 -1138
rect 581 -1144 584 -1138
rect 1252 -1145 1255 -1139
rect 1275 -1145 1278 -1139
rect 1306 -1145 1309 -1139
rect 1329 -1145 1332 -1139
rect 1407 -1144 1410 -1138
rect 1430 -1144 1433 -1138
rect 1461 -1144 1464 -1138
rect 1484 -1144 1487 -1138
rect 2120 -1144 2123 -1138
rect 2143 -1144 2146 -1138
rect 2174 -1144 2177 -1138
rect 2197 -1144 2200 -1138
rect 2275 -1143 2278 -1137
rect 2298 -1143 2301 -1137
rect 2329 -1143 2332 -1137
rect 2352 -1143 2355 -1137
rect -558 -1298 -555 -1292
rect -535 -1298 -532 -1292
rect -497 -1298 -494 -1292
rect -418 -1297 -415 -1291
rect -395 -1297 -392 -1291
rect -357 -1297 -354 -1291
rect -273 -1296 -270 -1290
rect -250 -1296 -247 -1290
rect -212 -1296 -209 -1290
rect -112 -1299 -109 -1293
rect -89 -1299 -86 -1293
rect -66 -1299 -63 -1293
rect -43 -1299 -40 -1293
rect 243 -1296 246 -1290
rect 266 -1296 269 -1290
rect 304 -1296 307 -1290
rect 383 -1295 386 -1289
rect 406 -1295 409 -1289
rect 444 -1295 447 -1289
rect 528 -1294 531 -1288
rect 551 -1294 554 -1288
rect 589 -1294 592 -1288
rect 689 -1297 692 -1291
rect 712 -1297 715 -1291
rect 735 -1297 738 -1291
rect 758 -1297 761 -1291
rect 1146 -1296 1149 -1290
rect 1169 -1296 1172 -1290
rect 1207 -1296 1210 -1290
rect 1286 -1295 1289 -1289
rect 1309 -1295 1312 -1289
rect 1347 -1295 1350 -1289
rect 1431 -1294 1434 -1288
rect 1454 -1294 1457 -1288
rect 1492 -1294 1495 -1288
rect 1592 -1297 1595 -1291
rect 1615 -1297 1618 -1291
rect 1638 -1297 1641 -1291
rect 1661 -1297 1664 -1291
rect 2014 -1295 2017 -1289
rect 2037 -1295 2040 -1289
rect 2075 -1295 2078 -1289
rect 2154 -1294 2157 -1288
rect 2177 -1294 2180 -1288
rect 2215 -1294 2218 -1288
rect 2299 -1293 2302 -1287
rect 2322 -1293 2325 -1287
rect 2360 -1293 2363 -1287
rect 2460 -1296 2463 -1290
rect 2483 -1296 2486 -1290
rect 2506 -1296 2509 -1290
rect 2529 -1296 2532 -1290
<< ndiffusion >>
rect -468 -889 -465 -885
rect -462 -889 -459 -885
rect -445 -889 -442 -885
rect -439 -889 -436 -885
rect -415 -889 -411 -885
rect -408 -889 -405 -885
rect -392 -889 -388 -885
rect -385 -889 -382 -885
rect 322 -889 325 -885
rect 328 -889 331 -885
rect 345 -889 348 -885
rect 351 -889 354 -885
rect 375 -889 379 -885
rect 382 -889 385 -885
rect 398 -889 402 -885
rect 405 -889 408 -885
rect 1304 -889 1307 -885
rect 1310 -889 1313 -885
rect 1327 -889 1330 -885
rect 1333 -889 1336 -885
rect 1357 -889 1361 -885
rect 1364 -889 1367 -885
rect 1380 -889 1384 -885
rect 1387 -889 1390 -885
rect 2188 -889 2191 -885
rect 2194 -889 2197 -885
rect 2211 -889 2214 -885
rect 2217 -889 2220 -885
rect 2241 -889 2245 -885
rect 2248 -889 2251 -885
rect 2264 -889 2268 -885
rect 2271 -889 2274 -885
rect -455 -1200 -452 -1196
rect -449 -1200 -446 -1196
rect -432 -1200 -429 -1196
rect -426 -1200 -423 -1196
rect -402 -1200 -398 -1196
rect -395 -1200 -392 -1196
rect -379 -1200 -375 -1196
rect -372 -1200 -369 -1196
rect -300 -1199 -297 -1195
rect -294 -1199 -291 -1195
rect -277 -1199 -274 -1195
rect -271 -1199 -268 -1195
rect -247 -1199 -243 -1195
rect -240 -1199 -237 -1195
rect -224 -1199 -220 -1195
rect -217 -1199 -214 -1195
rect 346 -1198 349 -1194
rect 352 -1198 355 -1194
rect 369 -1198 372 -1194
rect 375 -1198 378 -1194
rect 399 -1198 403 -1194
rect 406 -1198 409 -1194
rect 422 -1198 426 -1194
rect 429 -1198 432 -1194
rect 501 -1197 504 -1193
rect 507 -1197 510 -1193
rect 524 -1197 527 -1193
rect 530 -1197 533 -1193
rect 554 -1197 558 -1193
rect 561 -1197 564 -1193
rect 577 -1197 581 -1193
rect 584 -1197 587 -1193
rect 1249 -1198 1252 -1194
rect 1255 -1198 1258 -1194
rect 1272 -1198 1275 -1194
rect 1278 -1198 1281 -1194
rect 1302 -1198 1306 -1194
rect 1309 -1198 1312 -1194
rect 1325 -1198 1329 -1194
rect 1332 -1198 1335 -1194
rect 1404 -1197 1407 -1193
rect 1410 -1197 1413 -1193
rect 1427 -1197 1430 -1193
rect 1433 -1197 1436 -1193
rect 1457 -1197 1461 -1193
rect 1464 -1197 1467 -1193
rect 1480 -1197 1484 -1193
rect 1487 -1197 1490 -1193
rect 2117 -1197 2120 -1193
rect 2123 -1197 2126 -1193
rect 2140 -1197 2143 -1193
rect 2146 -1197 2149 -1193
rect 2170 -1197 2174 -1193
rect 2177 -1197 2180 -1193
rect 2193 -1197 2197 -1193
rect 2200 -1197 2203 -1193
rect 2272 -1196 2275 -1192
rect 2278 -1196 2281 -1192
rect 2295 -1196 2298 -1192
rect 2301 -1196 2304 -1192
rect 2325 -1196 2329 -1192
rect 2332 -1196 2335 -1192
rect 2348 -1196 2352 -1192
rect 2355 -1196 2358 -1192
rect -116 -1327 -112 -1322
rect -109 -1327 -106 -1322
rect -93 -1327 -89 -1322
rect -86 -1327 -83 -1322
rect -70 -1327 -66 -1322
rect -63 -1327 -60 -1322
rect -47 -1327 -43 -1322
rect -40 -1327 -37 -1322
rect 685 -1325 689 -1320
rect 692 -1325 695 -1320
rect 708 -1325 712 -1320
rect 715 -1325 718 -1320
rect 731 -1325 735 -1320
rect 738 -1325 741 -1320
rect 754 -1325 758 -1320
rect 761 -1325 764 -1320
rect -562 -1334 -558 -1329
rect -555 -1334 -552 -1329
rect -539 -1334 -535 -1329
rect -532 -1334 -529 -1329
rect -501 -1334 -497 -1329
rect -494 -1334 -491 -1329
rect -422 -1333 -418 -1328
rect -415 -1333 -412 -1328
rect -399 -1333 -395 -1328
rect -392 -1333 -389 -1328
rect -361 -1333 -357 -1328
rect -354 -1333 -351 -1328
rect -277 -1332 -273 -1327
rect -270 -1332 -267 -1327
rect -254 -1332 -250 -1327
rect -247 -1332 -244 -1327
rect -216 -1332 -212 -1327
rect -209 -1332 -206 -1327
rect 239 -1332 243 -1327
rect 246 -1332 249 -1327
rect 262 -1332 266 -1327
rect 269 -1332 272 -1327
rect 300 -1332 304 -1327
rect 307 -1332 310 -1327
rect 379 -1331 383 -1326
rect 386 -1331 389 -1326
rect 402 -1331 406 -1326
rect 409 -1331 412 -1326
rect 440 -1331 444 -1326
rect 447 -1331 450 -1326
rect 524 -1330 528 -1325
rect 531 -1330 534 -1325
rect 547 -1330 551 -1325
rect 554 -1330 557 -1325
rect 585 -1330 589 -1325
rect 592 -1330 595 -1325
rect 1588 -1325 1592 -1320
rect 1595 -1325 1598 -1320
rect 1611 -1325 1615 -1320
rect 1618 -1325 1621 -1320
rect 1634 -1325 1638 -1320
rect 1641 -1325 1644 -1320
rect 1657 -1325 1661 -1320
rect 1664 -1325 1667 -1320
rect 1142 -1332 1146 -1327
rect 1149 -1332 1152 -1327
rect 1165 -1332 1169 -1327
rect 1172 -1332 1175 -1327
rect 1203 -1332 1207 -1327
rect 1210 -1332 1213 -1327
rect 1282 -1331 1286 -1326
rect 1289 -1331 1292 -1326
rect 1305 -1331 1309 -1326
rect 1312 -1331 1315 -1326
rect 1343 -1331 1347 -1326
rect 1350 -1331 1353 -1326
rect 1427 -1330 1431 -1325
rect 1434 -1330 1437 -1325
rect 1450 -1330 1454 -1325
rect 1457 -1330 1460 -1325
rect 1488 -1330 1492 -1325
rect 1495 -1330 1498 -1325
rect 2456 -1324 2460 -1319
rect 2463 -1324 2466 -1319
rect 2479 -1324 2483 -1319
rect 2486 -1324 2489 -1319
rect 2502 -1324 2506 -1319
rect 2509 -1324 2512 -1319
rect 2525 -1324 2529 -1319
rect 2532 -1324 2535 -1319
rect 2010 -1331 2014 -1326
rect 2017 -1331 2020 -1326
rect 2033 -1331 2037 -1326
rect 2040 -1331 2043 -1326
rect 2071 -1331 2075 -1326
rect 2078 -1331 2081 -1326
rect 2150 -1330 2154 -1325
rect 2157 -1330 2160 -1325
rect 2173 -1330 2177 -1325
rect 2180 -1330 2183 -1325
rect 2211 -1330 2215 -1325
rect 2218 -1330 2221 -1325
rect 2295 -1329 2299 -1324
rect 2302 -1329 2305 -1324
rect 2318 -1329 2322 -1324
rect 2325 -1329 2328 -1324
rect 2356 -1329 2360 -1324
rect 2363 -1329 2366 -1324
<< pdiffusion >>
rect -468 -836 -465 -830
rect -462 -836 -459 -830
rect -445 -836 -442 -830
rect -439 -836 -436 -830
rect -414 -836 -411 -830
rect -408 -836 -405 -830
rect -391 -836 -388 -830
rect -385 -836 -382 -830
rect 322 -836 325 -830
rect 328 -836 331 -830
rect 345 -836 348 -830
rect 351 -836 354 -830
rect 376 -836 379 -830
rect 382 -836 385 -830
rect 399 -836 402 -830
rect 405 -836 408 -830
rect 1304 -836 1307 -830
rect 1310 -836 1313 -830
rect 1327 -836 1330 -830
rect 1333 -836 1336 -830
rect 1358 -836 1361 -830
rect 1364 -836 1367 -830
rect 1381 -836 1384 -830
rect 1387 -836 1390 -830
rect 2188 -836 2191 -830
rect 2194 -836 2197 -830
rect 2211 -836 2214 -830
rect 2217 -836 2220 -830
rect 2242 -836 2245 -830
rect 2248 -836 2251 -830
rect 2265 -836 2268 -830
rect 2271 -836 2274 -830
rect -455 -1147 -452 -1141
rect -449 -1147 -446 -1141
rect -432 -1147 -429 -1141
rect -426 -1147 -423 -1141
rect -401 -1147 -398 -1141
rect -395 -1147 -392 -1141
rect -378 -1147 -375 -1141
rect -372 -1147 -369 -1141
rect -300 -1146 -297 -1140
rect -294 -1146 -291 -1140
rect -277 -1146 -274 -1140
rect -271 -1146 -268 -1140
rect -246 -1146 -243 -1140
rect -240 -1146 -237 -1140
rect -223 -1146 -220 -1140
rect -217 -1146 -214 -1140
rect 346 -1145 349 -1139
rect 352 -1145 355 -1139
rect 369 -1145 372 -1139
rect 375 -1145 378 -1139
rect 400 -1145 403 -1139
rect 406 -1145 409 -1139
rect 423 -1145 426 -1139
rect 429 -1145 432 -1139
rect 501 -1144 504 -1138
rect 507 -1144 510 -1138
rect 524 -1144 527 -1138
rect 530 -1144 533 -1138
rect 555 -1144 558 -1138
rect 561 -1144 564 -1138
rect 578 -1144 581 -1138
rect 584 -1144 587 -1138
rect 1249 -1145 1252 -1139
rect 1255 -1145 1258 -1139
rect 1272 -1145 1275 -1139
rect 1278 -1145 1281 -1139
rect 1303 -1145 1306 -1139
rect 1309 -1145 1312 -1139
rect 1326 -1145 1329 -1139
rect 1332 -1145 1335 -1139
rect 1404 -1144 1407 -1138
rect 1410 -1144 1413 -1138
rect 1427 -1144 1430 -1138
rect 1433 -1144 1436 -1138
rect 1458 -1144 1461 -1138
rect 1464 -1144 1467 -1138
rect 1481 -1144 1484 -1138
rect 1487 -1144 1490 -1138
rect 2117 -1144 2120 -1138
rect 2123 -1144 2126 -1138
rect 2140 -1144 2143 -1138
rect 2146 -1144 2149 -1138
rect 2171 -1144 2174 -1138
rect 2177 -1144 2180 -1138
rect 2194 -1144 2197 -1138
rect 2200 -1144 2203 -1138
rect 2272 -1143 2275 -1137
rect 2278 -1143 2281 -1137
rect 2295 -1143 2298 -1137
rect 2301 -1143 2304 -1137
rect 2326 -1143 2329 -1137
rect 2332 -1143 2335 -1137
rect 2349 -1143 2352 -1137
rect 2355 -1143 2358 -1137
rect -561 -1298 -558 -1292
rect -555 -1298 -552 -1292
rect -538 -1298 -535 -1292
rect -532 -1298 -529 -1292
rect -500 -1298 -497 -1292
rect -494 -1298 -491 -1292
rect -421 -1297 -418 -1291
rect -415 -1297 -412 -1291
rect -398 -1297 -395 -1291
rect -392 -1297 -389 -1291
rect -360 -1297 -357 -1291
rect -354 -1297 -351 -1291
rect -276 -1296 -273 -1290
rect -270 -1296 -267 -1290
rect -253 -1296 -250 -1290
rect -247 -1296 -244 -1290
rect -215 -1296 -212 -1290
rect -209 -1296 -206 -1290
rect -115 -1299 -112 -1293
rect -109 -1299 -106 -1293
rect -92 -1299 -89 -1293
rect -86 -1299 -83 -1293
rect -69 -1299 -66 -1293
rect -63 -1299 -60 -1293
rect -46 -1299 -43 -1293
rect -40 -1299 -37 -1293
rect 240 -1296 243 -1290
rect 246 -1296 249 -1290
rect 263 -1296 266 -1290
rect 269 -1296 272 -1290
rect 301 -1296 304 -1290
rect 307 -1296 310 -1290
rect 380 -1295 383 -1289
rect 386 -1295 389 -1289
rect 403 -1295 406 -1289
rect 409 -1295 412 -1289
rect 441 -1295 444 -1289
rect 447 -1295 450 -1289
rect 525 -1294 528 -1288
rect 531 -1294 534 -1288
rect 548 -1294 551 -1288
rect 554 -1294 557 -1288
rect 586 -1294 589 -1288
rect 592 -1294 595 -1288
rect 686 -1297 689 -1291
rect 692 -1297 695 -1291
rect 709 -1297 712 -1291
rect 715 -1297 718 -1291
rect 732 -1297 735 -1291
rect 738 -1297 741 -1291
rect 755 -1297 758 -1291
rect 761 -1297 764 -1291
rect 1143 -1296 1146 -1290
rect 1149 -1296 1152 -1290
rect 1166 -1296 1169 -1290
rect 1172 -1296 1175 -1290
rect 1204 -1296 1207 -1290
rect 1210 -1296 1213 -1290
rect 1283 -1295 1286 -1289
rect 1289 -1295 1292 -1289
rect 1306 -1295 1309 -1289
rect 1312 -1295 1315 -1289
rect 1344 -1295 1347 -1289
rect 1350 -1295 1353 -1289
rect 1428 -1294 1431 -1288
rect 1434 -1294 1437 -1288
rect 1451 -1294 1454 -1288
rect 1457 -1294 1460 -1288
rect 1489 -1294 1492 -1288
rect 1495 -1294 1498 -1288
rect 1589 -1297 1592 -1291
rect 1595 -1297 1598 -1291
rect 1612 -1297 1615 -1291
rect 1618 -1297 1621 -1291
rect 1635 -1297 1638 -1291
rect 1641 -1297 1644 -1291
rect 1658 -1297 1661 -1291
rect 1664 -1297 1667 -1291
rect 2011 -1295 2014 -1289
rect 2017 -1295 2020 -1289
rect 2034 -1295 2037 -1289
rect 2040 -1295 2043 -1289
rect 2072 -1295 2075 -1289
rect 2078 -1295 2081 -1289
rect 2151 -1294 2154 -1288
rect 2157 -1294 2160 -1288
rect 2174 -1294 2177 -1288
rect 2180 -1294 2183 -1288
rect 2212 -1294 2215 -1288
rect 2218 -1294 2221 -1288
rect 2296 -1293 2299 -1287
rect 2302 -1293 2305 -1287
rect 2319 -1293 2322 -1287
rect 2325 -1293 2328 -1287
rect 2357 -1293 2360 -1287
rect 2363 -1293 2366 -1287
rect 2457 -1296 2460 -1290
rect 2463 -1296 2466 -1290
rect 2480 -1296 2483 -1290
rect 2486 -1296 2489 -1290
rect 2503 -1296 2506 -1290
rect 2509 -1296 2512 -1290
rect 2526 -1296 2529 -1290
rect 2532 -1296 2535 -1290
<< ndcontact >>
rect -473 -889 -468 -885
rect -459 -889 -455 -885
rect -450 -889 -445 -885
rect -436 -889 -432 -885
rect -419 -889 -415 -885
rect -405 -889 -401 -885
rect -396 -889 -392 -885
rect -382 -889 -378 -885
rect 317 -889 322 -885
rect 331 -889 335 -885
rect 340 -889 345 -885
rect 354 -889 358 -885
rect 371 -889 375 -885
rect 385 -889 389 -885
rect 394 -889 398 -885
rect 408 -889 412 -885
rect 1299 -889 1304 -885
rect 1313 -889 1317 -885
rect 1322 -889 1327 -885
rect 1336 -889 1340 -885
rect 1353 -889 1357 -885
rect 1367 -889 1371 -885
rect 1376 -889 1380 -885
rect 1390 -889 1394 -885
rect 2183 -889 2188 -885
rect 2197 -889 2201 -885
rect 2206 -889 2211 -885
rect 2220 -889 2224 -885
rect 2237 -889 2241 -885
rect 2251 -889 2255 -885
rect 2260 -889 2264 -885
rect 2274 -889 2278 -885
rect -460 -1200 -455 -1196
rect -446 -1200 -442 -1196
rect -437 -1200 -432 -1196
rect -423 -1200 -419 -1196
rect -406 -1200 -402 -1196
rect -392 -1200 -388 -1196
rect -383 -1200 -379 -1196
rect -369 -1200 -365 -1196
rect -305 -1199 -300 -1195
rect -291 -1199 -287 -1195
rect -282 -1199 -277 -1195
rect -268 -1199 -264 -1195
rect -251 -1199 -247 -1195
rect -237 -1199 -233 -1195
rect -228 -1199 -224 -1195
rect -214 -1199 -210 -1195
rect 341 -1198 346 -1194
rect 355 -1198 359 -1194
rect 364 -1198 369 -1194
rect 378 -1198 382 -1194
rect 395 -1198 399 -1194
rect 409 -1198 413 -1194
rect 418 -1198 422 -1194
rect 432 -1198 436 -1194
rect 496 -1197 501 -1193
rect 510 -1197 514 -1193
rect 519 -1197 524 -1193
rect 533 -1197 537 -1193
rect 550 -1197 554 -1193
rect 564 -1197 568 -1193
rect 573 -1197 577 -1193
rect 587 -1197 591 -1193
rect 1244 -1198 1249 -1194
rect 1258 -1198 1262 -1194
rect 1267 -1198 1272 -1194
rect 1281 -1198 1285 -1194
rect 1298 -1198 1302 -1194
rect 1312 -1198 1316 -1194
rect 1321 -1198 1325 -1194
rect 1335 -1198 1339 -1194
rect 1399 -1197 1404 -1193
rect 1413 -1197 1417 -1193
rect 1422 -1197 1427 -1193
rect 1436 -1197 1440 -1193
rect 1453 -1197 1457 -1193
rect 1467 -1197 1471 -1193
rect 1476 -1197 1480 -1193
rect 1490 -1197 1494 -1193
rect 2112 -1197 2117 -1193
rect 2126 -1197 2130 -1193
rect 2135 -1197 2140 -1193
rect 2149 -1197 2153 -1193
rect 2166 -1197 2170 -1193
rect 2180 -1197 2184 -1193
rect 2189 -1197 2193 -1193
rect 2203 -1197 2207 -1193
rect 2267 -1196 2272 -1192
rect 2281 -1196 2285 -1192
rect 2290 -1196 2295 -1192
rect 2304 -1196 2308 -1192
rect 2321 -1196 2325 -1192
rect 2335 -1196 2339 -1192
rect 2344 -1196 2348 -1192
rect 2358 -1196 2362 -1192
rect -120 -1327 -116 -1322
rect -106 -1327 -102 -1322
rect -97 -1327 -93 -1322
rect -83 -1327 -79 -1322
rect -74 -1327 -70 -1322
rect -60 -1327 -56 -1322
rect -51 -1327 -47 -1322
rect -37 -1327 -33 -1322
rect 681 -1325 685 -1320
rect 695 -1325 699 -1320
rect 704 -1325 708 -1320
rect 718 -1325 722 -1320
rect 727 -1325 731 -1320
rect 741 -1325 745 -1320
rect 750 -1325 754 -1320
rect 764 -1325 768 -1320
rect -566 -1334 -562 -1329
rect -552 -1334 -548 -1329
rect -543 -1334 -539 -1329
rect -529 -1334 -525 -1329
rect -505 -1334 -501 -1329
rect -491 -1334 -487 -1329
rect -426 -1333 -422 -1328
rect -412 -1333 -408 -1328
rect -403 -1333 -399 -1328
rect -389 -1333 -385 -1328
rect -365 -1333 -361 -1328
rect -351 -1333 -347 -1328
rect -281 -1332 -277 -1327
rect -267 -1332 -263 -1327
rect -258 -1332 -254 -1327
rect -244 -1332 -240 -1327
rect -220 -1332 -216 -1327
rect -206 -1332 -202 -1327
rect 235 -1332 239 -1327
rect 249 -1332 253 -1327
rect 258 -1332 262 -1327
rect 272 -1332 276 -1327
rect 296 -1332 300 -1327
rect 310 -1332 314 -1327
rect 375 -1331 379 -1326
rect 389 -1331 393 -1326
rect 398 -1331 402 -1326
rect 412 -1331 416 -1326
rect 436 -1331 440 -1326
rect 450 -1331 454 -1326
rect 520 -1330 524 -1325
rect 534 -1330 538 -1325
rect 543 -1330 547 -1325
rect 557 -1330 561 -1325
rect 581 -1330 585 -1325
rect 595 -1330 599 -1325
rect 1584 -1325 1588 -1320
rect 1598 -1325 1602 -1320
rect 1607 -1325 1611 -1320
rect 1621 -1325 1625 -1320
rect 1630 -1325 1634 -1320
rect 1644 -1325 1648 -1320
rect 1653 -1325 1657 -1320
rect 1667 -1325 1671 -1320
rect 1138 -1332 1142 -1327
rect 1152 -1332 1156 -1327
rect 1161 -1332 1165 -1327
rect 1175 -1332 1179 -1327
rect 1199 -1332 1203 -1327
rect 1213 -1332 1217 -1327
rect 1278 -1331 1282 -1326
rect 1292 -1331 1296 -1326
rect 1301 -1331 1305 -1326
rect 1315 -1331 1319 -1326
rect 1339 -1331 1343 -1326
rect 1353 -1331 1357 -1326
rect 1423 -1330 1427 -1325
rect 1437 -1330 1441 -1325
rect 1446 -1330 1450 -1325
rect 1460 -1330 1464 -1325
rect 1484 -1330 1488 -1325
rect 1498 -1330 1502 -1325
rect 2452 -1324 2456 -1319
rect 2466 -1324 2470 -1319
rect 2475 -1324 2479 -1319
rect 2489 -1324 2493 -1319
rect 2498 -1324 2502 -1319
rect 2512 -1324 2516 -1319
rect 2521 -1324 2525 -1319
rect 2535 -1324 2539 -1319
rect 2006 -1331 2010 -1326
rect 2020 -1331 2024 -1326
rect 2029 -1331 2033 -1326
rect 2043 -1331 2047 -1326
rect 2067 -1331 2071 -1326
rect 2081 -1331 2085 -1326
rect 2146 -1330 2150 -1325
rect 2160 -1330 2164 -1325
rect 2169 -1330 2173 -1325
rect 2183 -1330 2187 -1325
rect 2207 -1330 2211 -1325
rect 2221 -1330 2225 -1325
rect 2291 -1329 2295 -1324
rect 2305 -1329 2309 -1324
rect 2314 -1329 2318 -1324
rect 2328 -1329 2332 -1324
rect 2352 -1329 2356 -1324
rect 2366 -1329 2370 -1324
<< pdcontact >>
rect -473 -836 -468 -830
rect -459 -836 -455 -830
rect -450 -836 -445 -830
rect -436 -836 -432 -830
rect -419 -836 -414 -830
rect -405 -836 -401 -830
rect -396 -836 -391 -830
rect -382 -836 -378 -830
rect 317 -836 322 -830
rect 331 -836 335 -830
rect 340 -836 345 -830
rect 354 -836 358 -830
rect 371 -836 376 -830
rect 385 -836 389 -830
rect 394 -836 399 -830
rect 408 -836 412 -830
rect 1299 -836 1304 -830
rect 1313 -836 1317 -830
rect 1322 -836 1327 -830
rect 1336 -836 1340 -830
rect 1353 -836 1358 -830
rect 1367 -836 1371 -830
rect 1376 -836 1381 -830
rect 1390 -836 1394 -830
rect 2183 -836 2188 -830
rect 2197 -836 2201 -830
rect 2206 -836 2211 -830
rect 2220 -836 2224 -830
rect 2237 -836 2242 -830
rect 2251 -836 2255 -830
rect 2260 -836 2265 -830
rect 2274 -836 2278 -830
rect -460 -1147 -455 -1141
rect -446 -1147 -442 -1141
rect -437 -1147 -432 -1141
rect -423 -1147 -419 -1141
rect -406 -1147 -401 -1141
rect -392 -1147 -388 -1141
rect -383 -1147 -378 -1141
rect -369 -1147 -365 -1141
rect -305 -1146 -300 -1140
rect -291 -1146 -287 -1140
rect -282 -1146 -277 -1140
rect -268 -1146 -264 -1140
rect -251 -1146 -246 -1140
rect -237 -1146 -233 -1140
rect -228 -1146 -223 -1140
rect -214 -1146 -210 -1140
rect 341 -1145 346 -1139
rect 355 -1145 359 -1139
rect 364 -1145 369 -1139
rect 378 -1145 382 -1139
rect 395 -1145 400 -1139
rect 409 -1145 413 -1139
rect 418 -1145 423 -1139
rect 432 -1145 436 -1139
rect 496 -1144 501 -1138
rect 510 -1144 514 -1138
rect 519 -1144 524 -1138
rect 533 -1144 537 -1138
rect 550 -1144 555 -1138
rect 564 -1144 568 -1138
rect 573 -1144 578 -1138
rect 587 -1144 591 -1138
rect 1244 -1145 1249 -1139
rect 1258 -1145 1262 -1139
rect 1267 -1145 1272 -1139
rect 1281 -1145 1285 -1139
rect 1298 -1145 1303 -1139
rect 1312 -1145 1316 -1139
rect 1321 -1145 1326 -1139
rect 1335 -1145 1339 -1139
rect 1399 -1144 1404 -1138
rect 1413 -1144 1417 -1138
rect 1422 -1144 1427 -1138
rect 1436 -1144 1440 -1138
rect 1453 -1144 1458 -1138
rect 1467 -1144 1471 -1138
rect 1476 -1144 1481 -1138
rect 1490 -1144 1494 -1138
rect 2112 -1144 2117 -1138
rect 2126 -1144 2130 -1138
rect 2135 -1144 2140 -1138
rect 2149 -1144 2153 -1138
rect 2166 -1144 2171 -1138
rect 2180 -1144 2184 -1138
rect 2189 -1144 2194 -1138
rect 2203 -1144 2207 -1138
rect 2267 -1143 2272 -1137
rect 2281 -1143 2285 -1137
rect 2290 -1143 2295 -1137
rect 2304 -1143 2308 -1137
rect 2321 -1143 2326 -1137
rect 2335 -1143 2339 -1137
rect 2344 -1143 2349 -1137
rect 2358 -1143 2362 -1137
rect -566 -1298 -561 -1292
rect -552 -1298 -548 -1292
rect -543 -1298 -538 -1292
rect -529 -1298 -525 -1292
rect -505 -1298 -500 -1292
rect -491 -1298 -487 -1292
rect -426 -1297 -421 -1291
rect -412 -1297 -408 -1291
rect -403 -1297 -398 -1291
rect -389 -1297 -385 -1291
rect -365 -1297 -360 -1291
rect -351 -1297 -347 -1291
rect -281 -1296 -276 -1290
rect -267 -1296 -263 -1290
rect -258 -1296 -253 -1290
rect -244 -1296 -240 -1290
rect -220 -1296 -215 -1290
rect -206 -1296 -202 -1290
rect -120 -1299 -115 -1293
rect -106 -1299 -102 -1293
rect -97 -1299 -92 -1293
rect -83 -1299 -79 -1293
rect -74 -1299 -69 -1293
rect -60 -1299 -56 -1293
rect -51 -1299 -46 -1293
rect -37 -1299 -33 -1293
rect 235 -1296 240 -1290
rect 249 -1296 253 -1290
rect 258 -1296 263 -1290
rect 272 -1296 276 -1290
rect 296 -1296 301 -1290
rect 310 -1296 314 -1290
rect 375 -1295 380 -1289
rect 389 -1295 393 -1289
rect 398 -1295 403 -1289
rect 412 -1295 416 -1289
rect 436 -1295 441 -1289
rect 450 -1295 454 -1289
rect 520 -1294 525 -1288
rect 534 -1294 538 -1288
rect 543 -1294 548 -1288
rect 557 -1294 561 -1288
rect 581 -1294 586 -1288
rect 595 -1294 599 -1288
rect 681 -1297 686 -1291
rect 695 -1297 699 -1291
rect 704 -1297 709 -1291
rect 718 -1297 722 -1291
rect 727 -1297 732 -1291
rect 741 -1297 745 -1291
rect 750 -1297 755 -1291
rect 764 -1297 768 -1291
rect 1138 -1296 1143 -1290
rect 1152 -1296 1156 -1290
rect 1161 -1296 1166 -1290
rect 1175 -1296 1179 -1290
rect 1199 -1296 1204 -1290
rect 1213 -1296 1217 -1290
rect 1278 -1295 1283 -1289
rect 1292 -1295 1296 -1289
rect 1301 -1295 1306 -1289
rect 1315 -1295 1319 -1289
rect 1339 -1295 1344 -1289
rect 1353 -1295 1357 -1289
rect 1423 -1294 1428 -1288
rect 1437 -1294 1441 -1288
rect 1446 -1294 1451 -1288
rect 1460 -1294 1464 -1288
rect 1484 -1294 1489 -1288
rect 1498 -1294 1502 -1288
rect 1584 -1297 1589 -1291
rect 1598 -1297 1602 -1291
rect 1607 -1297 1612 -1291
rect 1621 -1297 1625 -1291
rect 1630 -1297 1635 -1291
rect 1644 -1297 1648 -1291
rect 1653 -1297 1658 -1291
rect 1667 -1297 1671 -1291
rect 2006 -1295 2011 -1289
rect 2020 -1295 2024 -1289
rect 2029 -1295 2034 -1289
rect 2043 -1295 2047 -1289
rect 2067 -1295 2072 -1289
rect 2081 -1295 2085 -1289
rect 2146 -1294 2151 -1288
rect 2160 -1294 2164 -1288
rect 2169 -1294 2174 -1288
rect 2183 -1294 2187 -1288
rect 2207 -1294 2212 -1288
rect 2221 -1294 2225 -1288
rect 2291 -1293 2296 -1287
rect 2305 -1293 2309 -1287
rect 2314 -1293 2319 -1287
rect 2328 -1293 2332 -1287
rect 2352 -1293 2357 -1287
rect 2366 -1293 2370 -1287
rect 2452 -1296 2457 -1290
rect 2466 -1296 2470 -1290
rect 2475 -1296 2480 -1290
rect 2489 -1296 2493 -1290
rect 2498 -1296 2503 -1290
rect 2512 -1296 2516 -1290
rect 2521 -1296 2526 -1290
rect 2535 -1296 2539 -1290
<< polysilicon >>
rect -489 -811 -439 -808
rect -489 -906 -486 -811
rect -465 -830 -462 -826
rect -442 -830 -439 -811
rect -411 -830 -408 -826
rect -388 -830 -385 -773
rect 301 -811 351 -808
rect -465 -875 -462 -836
rect -442 -842 -439 -836
rect -411 -854 -408 -836
rect -413 -858 -408 -854
rect -465 -878 -439 -875
rect -465 -885 -462 -881
rect -442 -885 -439 -878
rect -411 -885 -408 -858
rect -388 -885 -385 -836
rect -465 -906 -462 -889
rect -442 -893 -439 -889
rect -411 -892 -408 -889
rect -388 -891 -385 -889
rect -400 -893 -385 -891
rect -442 -895 -420 -893
rect -422 -897 -420 -895
rect -400 -897 -398 -893
rect -422 -899 -398 -897
rect -369 -906 -366 -858
rect -489 -909 -366 -906
rect 301 -906 304 -811
rect 325 -830 328 -826
rect 348 -830 351 -811
rect 379 -830 382 -826
rect 402 -830 405 -773
rect 1283 -811 1333 -808
rect 325 -875 328 -836
rect 348 -842 351 -836
rect 379 -854 382 -836
rect 377 -858 382 -854
rect 325 -878 351 -875
rect 325 -885 328 -881
rect 348 -885 351 -878
rect 379 -885 382 -858
rect 402 -885 405 -836
rect 325 -906 328 -889
rect 348 -893 351 -889
rect 379 -892 382 -889
rect 402 -891 405 -889
rect 390 -893 405 -891
rect 348 -895 370 -893
rect 368 -897 370 -895
rect 390 -897 392 -893
rect 368 -899 392 -897
rect 421 -906 424 -858
rect 301 -909 424 -906
rect 1283 -906 1286 -811
rect 1307 -830 1310 -826
rect 1330 -830 1333 -811
rect 1361 -830 1364 -826
rect 1384 -830 1387 -773
rect 2167 -811 2217 -808
rect 1307 -875 1310 -836
rect 1330 -842 1333 -836
rect 1361 -854 1364 -836
rect 1359 -858 1364 -854
rect 1307 -878 1333 -875
rect 1307 -885 1310 -881
rect 1330 -885 1333 -878
rect 1361 -885 1364 -858
rect 1384 -885 1387 -836
rect 1307 -906 1310 -889
rect 1330 -893 1333 -889
rect 1361 -892 1364 -889
rect 1384 -891 1387 -889
rect 1372 -893 1387 -891
rect 1330 -895 1352 -893
rect 1350 -897 1352 -895
rect 1372 -897 1374 -893
rect 1350 -899 1374 -897
rect 1403 -906 1406 -858
rect 1283 -909 1406 -906
rect 2167 -906 2170 -811
rect 2191 -830 2194 -826
rect 2214 -830 2217 -811
rect 2245 -830 2248 -826
rect 2268 -830 2271 -773
rect 2191 -875 2194 -836
rect 2214 -842 2217 -836
rect 2245 -854 2248 -836
rect 2243 -858 2248 -854
rect 2191 -878 2217 -875
rect 2191 -885 2194 -881
rect 2214 -885 2217 -878
rect 2245 -885 2248 -858
rect 2268 -885 2271 -836
rect 2191 -906 2194 -889
rect 2214 -893 2217 -889
rect 2245 -892 2248 -889
rect 2268 -891 2271 -889
rect 2256 -893 2271 -891
rect 2214 -895 2236 -893
rect 2234 -897 2236 -895
rect 2256 -897 2258 -893
rect 2234 -899 2258 -897
rect 2287 -906 2290 -858
rect 2167 -909 2290 -906
rect -476 -1122 -426 -1119
rect -476 -1217 -473 -1122
rect -452 -1141 -449 -1137
rect -429 -1141 -426 -1122
rect -398 -1141 -395 -1137
rect -375 -1141 -372 -1078
rect -321 -1121 -271 -1118
rect -452 -1186 -449 -1147
rect -429 -1153 -426 -1147
rect -398 -1165 -395 -1147
rect -400 -1169 -395 -1165
rect -452 -1189 -426 -1186
rect -452 -1196 -449 -1192
rect -429 -1196 -426 -1189
rect -398 -1196 -395 -1169
rect -375 -1196 -372 -1147
rect -452 -1217 -449 -1200
rect -429 -1204 -426 -1200
rect -398 -1203 -395 -1200
rect -375 -1202 -372 -1200
rect -387 -1203 -372 -1202
rect -387 -1204 -376 -1203
rect -429 -1206 -407 -1204
rect -409 -1208 -407 -1206
rect -387 -1208 -385 -1204
rect -409 -1210 -385 -1208
rect -356 -1217 -351 -1169
rect -476 -1220 -351 -1217
rect -321 -1216 -318 -1121
rect -297 -1140 -294 -1136
rect -274 -1140 -271 -1121
rect -243 -1140 -240 -1136
rect -220 -1140 -217 -1112
rect 325 -1120 375 -1117
rect -297 -1185 -294 -1146
rect -274 -1152 -271 -1146
rect -243 -1164 -240 -1146
rect -245 -1168 -240 -1164
rect -297 -1188 -271 -1185
rect -297 -1195 -294 -1191
rect -274 -1195 -271 -1188
rect -243 -1195 -240 -1168
rect -220 -1195 -217 -1146
rect -297 -1216 -294 -1199
rect -274 -1203 -271 -1199
rect -243 -1202 -240 -1199
rect -220 -1201 -217 -1199
rect -232 -1202 -217 -1201
rect -232 -1203 -221 -1202
rect -274 -1205 -252 -1203
rect -254 -1207 -252 -1205
rect -232 -1207 -230 -1203
rect -254 -1209 -230 -1207
rect -201 -1216 -196 -1168
rect -321 -1219 -196 -1216
rect 325 -1215 328 -1120
rect 349 -1139 352 -1135
rect 372 -1139 375 -1120
rect 403 -1139 406 -1135
rect 426 -1139 429 -1069
rect 480 -1119 530 -1116
rect 349 -1184 352 -1145
rect 372 -1151 375 -1145
rect 403 -1163 406 -1145
rect 401 -1167 406 -1163
rect 349 -1187 375 -1184
rect 349 -1194 352 -1190
rect 372 -1194 375 -1187
rect 403 -1194 406 -1167
rect 426 -1194 429 -1145
rect 349 -1215 352 -1198
rect 372 -1202 375 -1198
rect 403 -1201 406 -1198
rect 426 -1200 429 -1198
rect 414 -1201 429 -1200
rect 414 -1202 425 -1201
rect 372 -1204 394 -1202
rect 392 -1206 394 -1204
rect 414 -1206 416 -1202
rect 392 -1208 416 -1206
rect 445 -1215 450 -1167
rect 325 -1218 450 -1215
rect 480 -1214 483 -1119
rect 504 -1138 507 -1134
rect 527 -1138 530 -1119
rect 558 -1138 561 -1134
rect 581 -1138 584 -1116
rect 1228 -1120 1278 -1117
rect 504 -1183 507 -1144
rect 527 -1150 530 -1144
rect 558 -1162 561 -1144
rect 556 -1166 561 -1162
rect 504 -1186 530 -1183
rect 504 -1193 507 -1189
rect 527 -1193 530 -1186
rect 558 -1193 561 -1166
rect 581 -1193 584 -1144
rect 504 -1214 507 -1197
rect 527 -1201 530 -1197
rect 558 -1200 561 -1197
rect 581 -1199 584 -1197
rect 569 -1200 584 -1199
rect 569 -1201 580 -1200
rect 527 -1203 549 -1201
rect 547 -1205 549 -1203
rect 569 -1205 571 -1201
rect 547 -1207 571 -1205
rect 600 -1214 605 -1166
rect 480 -1217 605 -1214
rect 1228 -1215 1231 -1120
rect 1252 -1139 1255 -1135
rect 1275 -1139 1278 -1120
rect 1306 -1139 1309 -1135
rect 1329 -1139 1332 -1069
rect 1383 -1119 1433 -1116
rect 1252 -1184 1255 -1145
rect 1275 -1151 1278 -1145
rect 1306 -1163 1309 -1145
rect 1304 -1167 1309 -1163
rect 1252 -1187 1278 -1184
rect 1252 -1194 1255 -1190
rect 1275 -1194 1278 -1187
rect 1306 -1194 1309 -1167
rect 1329 -1194 1332 -1145
rect 1252 -1215 1255 -1198
rect 1275 -1202 1278 -1198
rect 1306 -1201 1309 -1198
rect 1329 -1200 1332 -1198
rect 1317 -1201 1332 -1200
rect 1317 -1202 1328 -1201
rect 1275 -1204 1297 -1202
rect 1295 -1206 1297 -1204
rect 1317 -1206 1319 -1202
rect 1295 -1208 1319 -1206
rect 1348 -1215 1353 -1167
rect 1228 -1218 1353 -1215
rect 1383 -1214 1386 -1119
rect 1407 -1138 1410 -1134
rect 1430 -1138 1433 -1119
rect 1461 -1138 1464 -1134
rect 1484 -1138 1487 -1118
rect 2096 -1119 2146 -1116
rect 1407 -1183 1410 -1144
rect 1430 -1150 1433 -1144
rect 1461 -1162 1464 -1144
rect 1459 -1166 1464 -1162
rect 1407 -1186 1433 -1183
rect 1407 -1193 1410 -1189
rect 1430 -1193 1433 -1186
rect 1461 -1193 1464 -1166
rect 1484 -1193 1487 -1144
rect 1407 -1214 1410 -1197
rect 1430 -1201 1433 -1197
rect 1461 -1200 1464 -1197
rect 1484 -1199 1487 -1197
rect 1472 -1200 1487 -1199
rect 1472 -1201 1483 -1200
rect 1430 -1203 1452 -1201
rect 1450 -1205 1452 -1203
rect 1472 -1205 1474 -1201
rect 1450 -1207 1474 -1205
rect 1503 -1214 1508 -1166
rect 1383 -1217 1508 -1214
rect 2096 -1214 2099 -1119
rect 2120 -1138 2123 -1134
rect 2143 -1138 2146 -1119
rect 2174 -1138 2177 -1134
rect 2197 -1138 2200 -1069
rect 2251 -1118 2301 -1115
rect 2120 -1183 2123 -1144
rect 2143 -1150 2146 -1144
rect 2174 -1162 2177 -1144
rect 2172 -1166 2177 -1162
rect 2120 -1186 2146 -1183
rect 2120 -1193 2123 -1189
rect 2143 -1193 2146 -1186
rect 2174 -1193 2177 -1166
rect 2197 -1193 2200 -1144
rect 2120 -1214 2123 -1197
rect 2143 -1201 2146 -1197
rect 2174 -1200 2177 -1197
rect 2197 -1199 2200 -1197
rect 2185 -1200 2200 -1199
rect 2185 -1201 2196 -1200
rect 2143 -1203 2165 -1201
rect 2163 -1205 2165 -1203
rect 2185 -1205 2187 -1201
rect 2163 -1207 2187 -1205
rect 2216 -1214 2221 -1166
rect 2096 -1217 2221 -1214
rect 2251 -1213 2254 -1118
rect 2275 -1137 2278 -1133
rect 2298 -1137 2301 -1118
rect 2329 -1137 2332 -1133
rect 2352 -1137 2355 -1118
rect 2275 -1182 2278 -1143
rect 2298 -1149 2301 -1143
rect 2329 -1161 2332 -1143
rect 2327 -1165 2332 -1161
rect 2275 -1185 2301 -1182
rect 2275 -1192 2278 -1188
rect 2298 -1192 2301 -1185
rect 2329 -1192 2332 -1165
rect 2352 -1192 2355 -1143
rect 2275 -1213 2278 -1196
rect 2298 -1200 2301 -1196
rect 2329 -1199 2332 -1196
rect 2352 -1198 2355 -1196
rect 2340 -1199 2355 -1198
rect 2340 -1200 2351 -1199
rect 2298 -1202 2320 -1200
rect 2318 -1204 2320 -1202
rect 2340 -1204 2342 -1200
rect 2318 -1206 2342 -1204
rect 2371 -1213 2376 -1165
rect 2251 -1216 2376 -1213
rect -558 -1292 -555 -1289
rect -535 -1292 -532 -1289
rect -497 -1292 -494 -1289
rect -418 -1291 -415 -1288
rect -395 -1291 -392 -1288
rect -357 -1291 -354 -1288
rect -273 -1290 -270 -1287
rect -250 -1290 -247 -1287
rect -212 -1290 -209 -1287
rect -112 -1293 -109 -1289
rect -89 -1293 -86 -1289
rect -66 -1293 -63 -1289
rect -43 -1293 -40 -1289
rect 243 -1290 246 -1287
rect 266 -1290 269 -1287
rect 304 -1290 307 -1287
rect 383 -1289 386 -1286
rect 406 -1289 409 -1286
rect 444 -1289 447 -1286
rect 528 -1288 531 -1285
rect 551 -1288 554 -1285
rect 589 -1288 592 -1285
rect -558 -1309 -555 -1298
rect -560 -1313 -555 -1309
rect -558 -1329 -555 -1313
rect -535 -1318 -532 -1298
rect -497 -1308 -494 -1298
rect -418 -1308 -415 -1297
rect -499 -1312 -494 -1308
rect -420 -1312 -415 -1308
rect -537 -1322 -532 -1318
rect -535 -1329 -532 -1322
rect -497 -1329 -494 -1312
rect -418 -1328 -415 -1312
rect -395 -1317 -392 -1297
rect -357 -1307 -354 -1297
rect -273 -1307 -270 -1296
rect -359 -1311 -354 -1307
rect -275 -1311 -270 -1307
rect -397 -1321 -392 -1317
rect -395 -1328 -392 -1321
rect -357 -1328 -354 -1311
rect -273 -1327 -270 -1311
rect -250 -1316 -247 -1296
rect -212 -1306 -209 -1296
rect 689 -1291 692 -1287
rect 712 -1291 715 -1287
rect 735 -1291 738 -1287
rect 758 -1291 761 -1287
rect 1146 -1290 1149 -1287
rect 1169 -1290 1172 -1287
rect 1207 -1290 1210 -1287
rect 1286 -1289 1289 -1286
rect 1309 -1289 1312 -1286
rect 1347 -1289 1350 -1286
rect 1431 -1288 1434 -1285
rect 1454 -1288 1457 -1285
rect 1492 -1288 1495 -1285
rect -214 -1310 -209 -1306
rect -252 -1320 -247 -1316
rect -250 -1327 -247 -1320
rect -212 -1327 -209 -1310
rect -112 -1322 -109 -1299
rect -89 -1322 -86 -1299
rect -66 -1322 -63 -1299
rect -43 -1311 -40 -1299
rect 243 -1307 246 -1296
rect 241 -1311 246 -1307
rect -45 -1315 -40 -1311
rect -43 -1322 -40 -1315
rect 243 -1327 246 -1311
rect 266 -1316 269 -1296
rect 304 -1306 307 -1296
rect 383 -1306 386 -1295
rect 302 -1310 307 -1306
rect 381 -1310 386 -1306
rect 264 -1320 269 -1316
rect 266 -1327 269 -1320
rect 304 -1327 307 -1310
rect 383 -1326 386 -1310
rect 406 -1315 409 -1295
rect 444 -1305 447 -1295
rect 528 -1305 531 -1294
rect 442 -1309 447 -1305
rect 526 -1309 531 -1305
rect 404 -1319 409 -1315
rect 406 -1326 409 -1319
rect 444 -1326 447 -1309
rect 528 -1325 531 -1309
rect 551 -1314 554 -1294
rect 589 -1304 592 -1294
rect 1592 -1291 1595 -1287
rect 1615 -1291 1618 -1287
rect 1638 -1291 1641 -1287
rect 1661 -1291 1664 -1287
rect 2014 -1289 2017 -1286
rect 2037 -1289 2040 -1286
rect 2075 -1289 2078 -1286
rect 2154 -1288 2157 -1285
rect 2177 -1288 2180 -1285
rect 2215 -1288 2218 -1285
rect 2299 -1287 2302 -1284
rect 2322 -1287 2325 -1284
rect 2360 -1287 2363 -1284
rect 587 -1308 592 -1304
rect 549 -1318 554 -1314
rect 551 -1325 554 -1318
rect 589 -1325 592 -1308
rect 689 -1320 692 -1297
rect 712 -1320 715 -1297
rect 735 -1320 738 -1297
rect 758 -1309 761 -1297
rect 1146 -1307 1149 -1296
rect 756 -1313 761 -1309
rect 1144 -1311 1149 -1307
rect 758 -1320 761 -1313
rect -112 -1331 -109 -1327
rect -558 -1338 -555 -1334
rect -535 -1338 -532 -1334
rect -497 -1338 -494 -1334
rect -418 -1337 -415 -1333
rect -395 -1337 -392 -1333
rect -357 -1337 -354 -1333
rect -273 -1336 -270 -1332
rect -250 -1336 -247 -1332
rect -212 -1336 -209 -1332
rect -89 -1343 -86 -1327
rect -66 -1352 -63 -1327
rect -43 -1331 -40 -1327
rect 689 -1329 692 -1325
rect 243 -1336 246 -1332
rect 266 -1336 269 -1332
rect 304 -1336 307 -1332
rect 383 -1335 386 -1331
rect 406 -1335 409 -1331
rect 444 -1335 447 -1331
rect 528 -1334 531 -1330
rect 551 -1334 554 -1330
rect 589 -1334 592 -1330
rect 712 -1341 715 -1325
rect 735 -1350 738 -1325
rect 758 -1329 761 -1325
rect 1146 -1327 1149 -1311
rect 1169 -1316 1172 -1296
rect 1207 -1306 1210 -1296
rect 1286 -1306 1289 -1295
rect 1205 -1310 1210 -1306
rect 1284 -1310 1289 -1306
rect 1167 -1320 1172 -1316
rect 1169 -1327 1172 -1320
rect 1207 -1327 1210 -1310
rect 1286 -1326 1289 -1310
rect 1309 -1315 1312 -1295
rect 1347 -1305 1350 -1295
rect 1431 -1305 1434 -1294
rect 1345 -1309 1350 -1305
rect 1429 -1309 1434 -1305
rect 1307 -1319 1312 -1315
rect 1309 -1326 1312 -1319
rect 1347 -1326 1350 -1309
rect 1431 -1325 1434 -1309
rect 1454 -1314 1457 -1294
rect 1492 -1304 1495 -1294
rect 2460 -1290 2463 -1286
rect 2483 -1290 2486 -1286
rect 2506 -1290 2509 -1286
rect 2529 -1290 2532 -1286
rect 1490 -1308 1495 -1304
rect 1452 -1318 1457 -1314
rect 1454 -1325 1457 -1318
rect 1492 -1325 1495 -1308
rect 1592 -1320 1595 -1297
rect 1615 -1320 1618 -1297
rect 1638 -1320 1641 -1297
rect 1661 -1309 1664 -1297
rect 2014 -1306 2017 -1295
rect 1659 -1313 1664 -1309
rect 2012 -1310 2017 -1306
rect 1661 -1320 1664 -1313
rect 1592 -1329 1595 -1325
rect 1146 -1336 1149 -1332
rect 1169 -1336 1172 -1332
rect 1207 -1336 1210 -1332
rect 1286 -1335 1289 -1331
rect 1309 -1335 1312 -1331
rect 1347 -1335 1350 -1331
rect 1431 -1334 1434 -1330
rect 1454 -1334 1457 -1330
rect 1492 -1334 1495 -1330
rect 1615 -1341 1618 -1325
rect 1638 -1350 1641 -1325
rect 1661 -1329 1664 -1325
rect 2014 -1326 2017 -1310
rect 2037 -1315 2040 -1295
rect 2075 -1305 2078 -1295
rect 2154 -1305 2157 -1294
rect 2073 -1309 2078 -1305
rect 2152 -1309 2157 -1305
rect 2035 -1319 2040 -1315
rect 2037 -1326 2040 -1319
rect 2075 -1326 2078 -1309
rect 2154 -1325 2157 -1309
rect 2177 -1314 2180 -1294
rect 2215 -1304 2218 -1294
rect 2299 -1304 2302 -1293
rect 2213 -1308 2218 -1304
rect 2297 -1308 2302 -1304
rect 2175 -1318 2180 -1314
rect 2177 -1325 2180 -1318
rect 2215 -1325 2218 -1308
rect 2299 -1324 2302 -1308
rect 2322 -1313 2325 -1293
rect 2360 -1303 2363 -1293
rect 2358 -1307 2363 -1303
rect 2320 -1317 2325 -1313
rect 2322 -1324 2325 -1317
rect 2360 -1324 2363 -1307
rect 2460 -1319 2463 -1296
rect 2483 -1319 2486 -1296
rect 2506 -1319 2509 -1296
rect 2529 -1308 2532 -1296
rect 2527 -1312 2532 -1308
rect 2529 -1319 2532 -1312
rect 2460 -1328 2463 -1324
rect 2014 -1335 2017 -1331
rect 2037 -1335 2040 -1331
rect 2075 -1335 2078 -1331
rect 2154 -1334 2157 -1330
rect 2177 -1334 2180 -1330
rect 2215 -1334 2218 -1330
rect 2299 -1333 2302 -1329
rect 2322 -1333 2325 -1329
rect 2360 -1333 2363 -1329
rect 2483 -1340 2486 -1324
rect 2506 -1349 2509 -1324
rect 2529 -1328 2532 -1324
<< polycontact >>
rect -390 -773 -383 -768
rect 399 -773 406 -768
rect 1382 -773 1389 -768
rect 2268 -773 2272 -768
rect -418 -858 -413 -854
rect -369 -858 -365 -853
rect 372 -858 377 -854
rect 421 -858 425 -853
rect 1354 -858 1359 -854
rect 1403 -858 1407 -853
rect 2238 -858 2243 -854
rect 2287 -858 2291 -853
rect -379 -1078 -368 -1068
rect 423 -1069 431 -1062
rect 1327 -1069 1336 -1062
rect 2196 -1069 2205 -1062
rect -220 -1112 -214 -1104
rect -405 -1169 -400 -1165
rect -356 -1169 -351 -1165
rect -376 -1207 -371 -1203
rect -250 -1168 -245 -1164
rect -201 -1168 -196 -1164
rect -221 -1206 -216 -1202
rect 581 -1116 586 -1109
rect 396 -1167 401 -1163
rect 445 -1167 450 -1163
rect 425 -1205 430 -1201
rect 551 -1166 556 -1162
rect 600 -1166 605 -1162
rect 580 -1204 585 -1200
rect 1299 -1167 1304 -1163
rect 1348 -1167 1353 -1163
rect 1328 -1205 1333 -1201
rect 1484 -1118 1489 -1112
rect 1454 -1166 1459 -1162
rect 1503 -1166 1508 -1162
rect 1483 -1204 1488 -1200
rect 2167 -1166 2172 -1162
rect 2216 -1166 2221 -1162
rect 2196 -1204 2201 -1200
rect 2352 -1118 2358 -1113
rect 2322 -1165 2327 -1161
rect 2371 -1165 2376 -1161
rect 2351 -1203 2356 -1199
rect -565 -1313 -560 -1309
rect -504 -1312 -499 -1308
rect -425 -1312 -420 -1308
rect -542 -1322 -537 -1318
rect -364 -1311 -359 -1307
rect -280 -1311 -275 -1307
rect -402 -1321 -397 -1317
rect -219 -1310 -214 -1306
rect -117 -1310 -112 -1306
rect -257 -1320 -252 -1316
rect 236 -1311 241 -1307
rect -50 -1315 -45 -1311
rect 297 -1310 302 -1306
rect 376 -1310 381 -1306
rect 259 -1320 264 -1316
rect 437 -1309 442 -1305
rect 521 -1309 526 -1305
rect 399 -1319 404 -1315
rect 582 -1308 587 -1304
rect 684 -1308 689 -1304
rect 544 -1318 549 -1314
rect 751 -1313 756 -1309
rect 1139 -1311 1144 -1307
rect -89 -1347 -84 -1343
rect 712 -1345 717 -1341
rect 1200 -1310 1205 -1306
rect 1279 -1310 1284 -1306
rect 1162 -1320 1167 -1316
rect 1340 -1309 1345 -1305
rect 1424 -1309 1429 -1305
rect 1302 -1319 1307 -1315
rect 1485 -1308 1490 -1304
rect 1587 -1308 1592 -1304
rect 1447 -1318 1452 -1314
rect 1654 -1313 1659 -1309
rect 2007 -1310 2012 -1306
rect 1615 -1345 1620 -1341
rect 2068 -1309 2073 -1305
rect 2147 -1309 2152 -1305
rect 2030 -1319 2035 -1315
rect 2208 -1308 2213 -1304
rect 2292 -1308 2297 -1304
rect 2170 -1318 2175 -1314
rect 2353 -1307 2358 -1303
rect 2455 -1307 2460 -1303
rect 2315 -1317 2320 -1313
rect 2522 -1312 2527 -1308
rect 2483 -1344 2488 -1340
rect -67 -1356 -62 -1352
rect 734 -1354 739 -1350
rect 1637 -1354 1642 -1350
rect 2505 -1353 2510 -1349
<< metal1 >>
rect -771 -933 -762 -770
rect -722 -782 -713 -770
rect -392 -773 -390 -768
rect -383 -773 399 -768
rect 406 -773 1382 -768
rect 1389 -773 2268 -768
rect 2272 -772 2389 -768
rect -722 -789 2281 -782
rect -771 -1341 -762 -943
rect -722 -1102 -713 -789
rect -473 -805 -424 -801
rect -473 -830 -468 -805
rect -473 -885 -468 -836
rect -459 -820 -432 -815
rect -459 -830 -455 -820
rect -436 -830 -432 -820
rect -459 -885 -455 -836
rect -459 -924 -455 -889
rect -450 -885 -445 -836
rect -436 -885 -432 -836
rect -427 -854 -424 -805
rect -419 -813 -415 -789
rect 317 -805 366 -801
rect -419 -818 -391 -813
rect -419 -830 -414 -818
rect -396 -830 -391 -818
rect 317 -830 322 -805
rect -427 -858 -418 -854
rect -405 -863 -401 -836
rect -427 -867 -401 -863
rect -450 -897 -445 -889
rect -427 -897 -424 -867
rect -405 -885 -401 -867
rect -382 -853 -378 -836
rect -382 -858 -369 -853
rect -382 -885 -378 -858
rect -450 -900 -424 -897
rect 317 -885 322 -836
rect 331 -820 358 -815
rect 331 -830 335 -820
rect 354 -830 358 -820
rect 331 -885 335 -836
rect -419 -900 -415 -889
rect -396 -900 -392 -889
rect -419 -904 -392 -900
rect -419 -933 -415 -904
rect 331 -924 335 -889
rect 340 -885 345 -836
rect 354 -885 358 -836
rect 363 -854 366 -805
rect 371 -813 375 -789
rect 1299 -805 1348 -801
rect 371 -818 399 -813
rect 371 -830 376 -818
rect 394 -830 399 -818
rect 1299 -830 1304 -805
rect 363 -858 372 -854
rect 385 -863 389 -836
rect 363 -867 389 -863
rect 340 -897 345 -889
rect 363 -897 366 -867
rect 385 -885 389 -867
rect 408 -853 412 -836
rect 408 -858 421 -853
rect 408 -885 412 -858
rect 340 -900 366 -897
rect 1299 -885 1304 -836
rect 1313 -820 1340 -815
rect 1313 -830 1317 -820
rect 1336 -830 1340 -820
rect 1313 -885 1317 -836
rect 371 -900 375 -889
rect 394 -900 398 -889
rect 371 -904 398 -900
rect 371 -932 375 -904
rect 1313 -924 1317 -889
rect 1322 -885 1327 -836
rect 1336 -885 1340 -836
rect 1345 -854 1348 -805
rect 1353 -813 1357 -789
rect 2183 -805 2232 -801
rect 1353 -818 1381 -813
rect 1353 -830 1358 -818
rect 1376 -830 1381 -818
rect 2183 -830 2188 -805
rect 1345 -858 1354 -854
rect 1367 -863 1371 -836
rect 1345 -867 1371 -863
rect 1322 -897 1327 -889
rect 1345 -897 1348 -867
rect 1367 -885 1371 -867
rect 1390 -853 1394 -836
rect 1390 -858 1403 -853
rect 1390 -885 1394 -858
rect 1322 -900 1348 -897
rect 2183 -885 2188 -836
rect 2197 -820 2224 -815
rect 2197 -830 2201 -820
rect 2220 -830 2224 -820
rect 2197 -885 2201 -836
rect 1353 -900 1357 -889
rect 1376 -900 1380 -889
rect 1353 -904 1380 -900
rect 1353 -932 1357 -904
rect 2197 -923 2201 -889
rect 2206 -885 2211 -836
rect 2220 -885 2224 -836
rect 2229 -854 2232 -805
rect 2237 -813 2241 -789
rect 2237 -818 2265 -813
rect 2237 -830 2242 -818
rect 2260 -830 2265 -818
rect 2229 -858 2238 -854
rect 2251 -863 2255 -836
rect 2229 -867 2255 -863
rect 2206 -897 2211 -889
rect 2229 -897 2232 -867
rect 2251 -885 2255 -867
rect 2274 -853 2278 -836
rect 2274 -858 2287 -853
rect 2274 -885 2278 -858
rect 2206 -900 2232 -897
rect 2237 -900 2241 -889
rect 2260 -900 2264 -889
rect 2237 -904 2264 -900
rect 2237 -932 2241 -904
rect -196 -933 2288 -932
rect -676 -940 2288 -933
rect -460 -1071 -455 -957
rect 330 -1063 335 -949
rect 330 -1068 423 -1063
rect -460 -1078 -379 -1071
rect 1313 -1063 1318 -948
rect 2197 -1062 2202 -952
rect 1313 -1069 1327 -1063
rect -244 -1090 2377 -1080
rect -243 -1102 -237 -1090
rect 558 -1100 564 -1090
rect 1461 -1100 1467 -1090
rect 2329 -1100 2335 -1090
rect -722 -1107 -237 -1102
rect 50 -1104 63 -1103
rect -678 -1270 -673 -1107
rect -460 -1116 -411 -1112
rect -460 -1141 -455 -1116
rect -654 -1237 -508 -1233
rect -654 -1341 -648 -1237
rect -493 -1250 -490 -1170
rect -460 -1196 -455 -1147
rect -446 -1131 -424 -1126
rect -446 -1141 -442 -1131
rect -423 -1141 -419 -1131
rect -446 -1196 -442 -1147
rect -437 -1196 -432 -1147
rect -423 -1196 -419 -1147
rect -414 -1165 -411 -1116
rect -399 -1124 -396 -1107
rect -300 -1115 -256 -1111
rect -406 -1129 -378 -1124
rect -406 -1141 -401 -1129
rect -383 -1141 -378 -1129
rect -305 -1140 -300 -1116
rect -411 -1169 -405 -1165
rect -392 -1174 -388 -1147
rect -414 -1178 -388 -1174
rect -437 -1208 -432 -1200
rect -414 -1208 -411 -1178
rect -392 -1196 -388 -1178
rect -369 -1165 -365 -1147
rect -369 -1169 -356 -1165
rect -369 -1196 -365 -1169
rect -437 -1211 -411 -1208
rect -305 -1195 -300 -1146
rect -291 -1130 -264 -1125
rect -291 -1140 -287 -1130
rect -268 -1140 -264 -1130
rect -291 -1195 -287 -1146
rect -282 -1195 -277 -1146
rect -268 -1195 -264 -1146
rect -259 -1164 -256 -1115
rect -240 -1123 -237 -1107
rect -214 -1112 63 -1104
rect -251 -1128 -223 -1123
rect -251 -1140 -246 -1128
rect -228 -1140 -223 -1128
rect -259 -1168 -250 -1164
rect -237 -1173 -233 -1146
rect -259 -1177 -233 -1173
rect -406 -1211 -402 -1200
rect -383 -1211 -379 -1200
rect -282 -1207 -277 -1199
rect -259 -1207 -256 -1177
rect -237 -1195 -233 -1177
rect -214 -1164 -210 -1146
rect -214 -1168 -201 -1164
rect -214 -1195 -210 -1168
rect -406 -1215 -379 -1211
rect -394 -1233 -391 -1215
rect -375 -1221 -372 -1207
rect -282 -1210 -256 -1207
rect -251 -1210 -247 -1199
rect -228 -1210 -224 -1199
rect -251 -1214 -224 -1210
rect -237 -1233 -234 -1214
rect -461 -1237 -234 -1233
rect -220 -1242 -217 -1206
rect -441 -1246 -217 -1242
rect -606 -1254 -322 -1250
rect -606 -1309 -600 -1254
rect -589 -1261 -584 -1260
rect -589 -1264 -376 -1261
rect -589 -1265 -584 -1264
rect -588 -1297 -585 -1265
rect -541 -1282 -538 -1275
rect -573 -1286 -479 -1282
rect -566 -1292 -561 -1286
rect -543 -1292 -538 -1286
rect -505 -1292 -500 -1286
rect -552 -1308 -548 -1298
rect -529 -1308 -525 -1298
rect -491 -1308 -487 -1298
rect -606 -1313 -565 -1309
rect -552 -1312 -504 -1308
rect -491 -1312 -478 -1308
rect -584 -1322 -542 -1318
rect -529 -1329 -525 -1312
rect -491 -1329 -487 -1312
rect -771 -1343 -648 -1341
rect -548 -1334 -543 -1329
rect -566 -1343 -562 -1334
rect -505 -1343 -501 -1334
rect -773 -1346 -505 -1343
rect -773 -1352 -648 -1346
rect -773 -1465 -758 -1352
rect -481 -1364 -478 -1312
rect -468 -1317 -463 -1264
rect -445 -1308 -442 -1272
rect -410 -1281 -407 -1275
rect -433 -1285 -339 -1281
rect -426 -1291 -421 -1285
rect -403 -1291 -398 -1285
rect -365 -1291 -360 -1285
rect -412 -1307 -408 -1297
rect -389 -1307 -385 -1297
rect -351 -1307 -347 -1297
rect -445 -1312 -425 -1308
rect -412 -1311 -364 -1307
rect -351 -1311 -340 -1307
rect -468 -1321 -402 -1317
rect -389 -1328 -385 -1311
rect -351 -1328 -347 -1311
rect -408 -1333 -403 -1328
rect -426 -1342 -422 -1333
rect -365 -1341 -361 -1333
rect -426 -1343 -365 -1342
rect -422 -1345 -365 -1343
rect -343 -1352 -340 -1311
rect -329 -1316 -322 -1254
rect -307 -1307 -301 -1246
rect -264 -1274 -101 -1271
rect -268 -1280 -265 -1275
rect -288 -1284 -194 -1280
rect -106 -1281 -101 -1274
rect -281 -1290 -276 -1284
rect -258 -1290 -253 -1284
rect -220 -1290 -215 -1284
rect -120 -1285 -46 -1281
rect -267 -1306 -263 -1296
rect -244 -1306 -240 -1296
rect -206 -1306 -202 -1296
rect -120 -1293 -115 -1285
rect -51 -1293 -46 -1285
rect -102 -1299 -97 -1293
rect -79 -1299 -74 -1293
rect -307 -1311 -280 -1307
rect -267 -1310 -219 -1306
rect -206 -1310 -117 -1306
rect -329 -1320 -257 -1316
rect -244 -1327 -240 -1310
rect -206 -1327 -202 -1310
rect -60 -1311 -56 -1299
rect -37 -1311 -33 -1299
rect -60 -1315 -50 -1311
rect -37 -1315 -28 -1311
rect -60 -1316 -56 -1315
rect -106 -1319 -56 -1316
rect -106 -1322 -102 -1319
rect -83 -1322 -79 -1319
rect -60 -1322 -56 -1319
rect -37 -1322 -33 -1315
rect -263 -1332 -258 -1327
rect -281 -1340 -277 -1332
rect -220 -1340 -216 -1332
rect -120 -1334 -116 -1327
rect -97 -1334 -93 -1327
rect -74 -1334 -70 -1327
rect -51 -1334 -47 -1327
rect -120 -1335 -47 -1334
rect -200 -1338 -47 -1335
rect -200 -1340 -195 -1338
rect -220 -1341 -195 -1340
rect -277 -1344 -195 -1341
rect -191 -1347 -89 -1344
rect -191 -1352 -187 -1347
rect -343 -1356 -187 -1352
rect -178 -1356 -67 -1352
rect -178 -1364 -175 -1356
rect -481 -1369 -175 -1364
rect 50 -1408 63 -1112
rect 123 -1105 564 -1100
rect 123 -1268 128 -1105
rect 341 -1114 390 -1110
rect 341 -1139 346 -1114
rect 147 -1235 293 -1231
rect 147 -1337 153 -1235
rect 308 -1248 311 -1168
rect 341 -1194 346 -1145
rect 355 -1129 377 -1124
rect 355 -1139 359 -1129
rect 378 -1139 382 -1129
rect 355 -1194 359 -1145
rect 364 -1194 369 -1145
rect 378 -1194 382 -1145
rect 387 -1163 390 -1114
rect 402 -1122 405 -1105
rect 501 -1113 545 -1109
rect 395 -1127 423 -1122
rect 395 -1139 400 -1127
rect 418 -1139 423 -1127
rect 496 -1138 501 -1114
rect 390 -1167 396 -1163
rect 409 -1172 413 -1145
rect 387 -1176 413 -1172
rect 364 -1206 369 -1198
rect 387 -1206 390 -1176
rect 409 -1194 413 -1176
rect 432 -1163 436 -1145
rect 432 -1167 445 -1163
rect 432 -1194 436 -1167
rect 364 -1209 390 -1206
rect 496 -1193 501 -1144
rect 510 -1128 537 -1123
rect 510 -1138 514 -1128
rect 533 -1138 537 -1128
rect 510 -1193 514 -1144
rect 519 -1193 524 -1144
rect 533 -1193 537 -1144
rect 542 -1162 545 -1113
rect 561 -1121 564 -1105
rect 1026 -1105 1467 -1100
rect 586 -1116 892 -1109
rect 550 -1126 578 -1121
rect 550 -1138 555 -1126
rect 573 -1138 578 -1126
rect 542 -1166 551 -1162
rect 564 -1171 568 -1144
rect 542 -1175 568 -1171
rect 395 -1209 399 -1198
rect 418 -1209 422 -1198
rect 519 -1205 524 -1197
rect 542 -1205 545 -1175
rect 564 -1193 568 -1175
rect 587 -1162 591 -1144
rect 587 -1166 600 -1162
rect 587 -1193 591 -1166
rect 395 -1213 422 -1209
rect 407 -1231 410 -1213
rect 426 -1219 429 -1205
rect 519 -1208 545 -1205
rect 550 -1208 554 -1197
rect 573 -1208 577 -1197
rect 550 -1212 577 -1208
rect 564 -1231 567 -1212
rect 340 -1235 567 -1231
rect 581 -1240 584 -1204
rect 360 -1244 584 -1240
rect 195 -1252 479 -1248
rect 195 -1307 201 -1252
rect 212 -1259 217 -1258
rect 212 -1262 425 -1259
rect 212 -1263 217 -1262
rect 213 -1295 216 -1263
rect 260 -1280 263 -1273
rect 228 -1284 322 -1280
rect 235 -1290 240 -1284
rect 258 -1290 263 -1284
rect 296 -1290 301 -1284
rect 249 -1306 253 -1296
rect 272 -1306 276 -1296
rect 310 -1306 314 -1296
rect 195 -1311 236 -1307
rect 249 -1310 297 -1306
rect 310 -1310 323 -1306
rect 217 -1320 259 -1316
rect 272 -1327 276 -1310
rect 310 -1327 314 -1310
rect 253 -1332 258 -1327
rect 235 -1341 239 -1332
rect 296 -1341 300 -1332
rect 156 -1344 296 -1341
rect 320 -1362 323 -1310
rect 333 -1315 338 -1262
rect 356 -1306 359 -1270
rect 391 -1279 394 -1273
rect 368 -1283 462 -1279
rect 375 -1289 380 -1283
rect 398 -1289 403 -1283
rect 436 -1289 441 -1283
rect 389 -1305 393 -1295
rect 412 -1305 416 -1295
rect 450 -1305 454 -1295
rect 356 -1310 376 -1306
rect 389 -1309 437 -1305
rect 450 -1309 461 -1305
rect 333 -1319 399 -1315
rect 412 -1326 416 -1309
rect 450 -1326 454 -1309
rect 393 -1331 398 -1326
rect 375 -1340 379 -1331
rect 436 -1339 440 -1331
rect 375 -1341 436 -1340
rect 379 -1343 436 -1341
rect 458 -1350 461 -1309
rect 472 -1314 479 -1252
rect 494 -1305 500 -1244
rect 537 -1272 700 -1269
rect 533 -1278 536 -1273
rect 513 -1282 607 -1278
rect 695 -1279 700 -1272
rect 520 -1288 525 -1282
rect 543 -1288 548 -1282
rect 581 -1288 586 -1282
rect 681 -1283 755 -1279
rect 534 -1304 538 -1294
rect 557 -1304 561 -1294
rect 595 -1304 599 -1294
rect 681 -1291 686 -1283
rect 750 -1291 755 -1283
rect 699 -1297 704 -1291
rect 722 -1297 727 -1291
rect 494 -1309 521 -1305
rect 534 -1308 582 -1304
rect 595 -1308 684 -1304
rect 472 -1318 544 -1314
rect 557 -1325 561 -1308
rect 595 -1325 599 -1308
rect 741 -1309 745 -1297
rect 764 -1309 768 -1297
rect 741 -1313 751 -1309
rect 764 -1313 779 -1309
rect 741 -1314 745 -1313
rect 695 -1317 745 -1314
rect 695 -1320 699 -1317
rect 718 -1320 722 -1317
rect 741 -1320 745 -1317
rect 764 -1320 768 -1313
rect 538 -1330 543 -1325
rect 520 -1338 524 -1330
rect 581 -1338 585 -1330
rect 681 -1332 685 -1325
rect 704 -1332 708 -1325
rect 727 -1332 731 -1325
rect 750 -1332 754 -1325
rect 681 -1333 754 -1332
rect 601 -1336 754 -1333
rect 601 -1338 606 -1336
rect 581 -1339 606 -1338
rect 524 -1342 606 -1339
rect 610 -1345 712 -1342
rect 610 -1350 614 -1345
rect 458 -1354 614 -1350
rect 623 -1354 734 -1350
rect 623 -1362 626 -1354
rect 320 -1367 626 -1362
rect 772 -1408 779 -1313
rect 50 -1421 779 -1408
rect 878 -1403 892 -1116
rect 1026 -1268 1031 -1105
rect 1244 -1114 1293 -1110
rect 1244 -1139 1249 -1114
rect 1050 -1235 1196 -1231
rect 1050 -1340 1056 -1235
rect 1211 -1248 1214 -1168
rect 1244 -1194 1249 -1145
rect 1258 -1129 1280 -1124
rect 1258 -1139 1262 -1129
rect 1281 -1139 1285 -1129
rect 1258 -1194 1262 -1145
rect 1267 -1194 1272 -1145
rect 1281 -1194 1285 -1145
rect 1290 -1163 1293 -1114
rect 1305 -1122 1308 -1105
rect 1404 -1113 1448 -1109
rect 1298 -1127 1326 -1122
rect 1298 -1139 1303 -1127
rect 1321 -1139 1326 -1127
rect 1399 -1138 1404 -1114
rect 1293 -1167 1299 -1163
rect 1312 -1172 1316 -1145
rect 1290 -1176 1316 -1172
rect 1267 -1206 1272 -1198
rect 1290 -1206 1293 -1176
rect 1312 -1194 1316 -1176
rect 1335 -1163 1339 -1145
rect 1335 -1167 1348 -1163
rect 1335 -1194 1339 -1167
rect 1267 -1209 1293 -1206
rect 1399 -1193 1404 -1144
rect 1413 -1128 1440 -1123
rect 1413 -1138 1417 -1128
rect 1436 -1138 1440 -1128
rect 1413 -1193 1417 -1144
rect 1422 -1193 1427 -1144
rect 1436 -1193 1440 -1144
rect 1445 -1162 1448 -1113
rect 1464 -1121 1467 -1105
rect 1894 -1104 2335 -1100
rect 1719 -1112 1722 -1111
rect 1489 -1118 1722 -1112
rect 1453 -1126 1481 -1121
rect 1453 -1138 1458 -1126
rect 1476 -1138 1481 -1126
rect 1445 -1166 1454 -1162
rect 1467 -1171 1471 -1144
rect 1445 -1175 1471 -1171
rect 1298 -1209 1302 -1198
rect 1321 -1209 1325 -1198
rect 1422 -1205 1427 -1197
rect 1445 -1205 1448 -1175
rect 1467 -1193 1471 -1175
rect 1490 -1162 1494 -1144
rect 1490 -1166 1503 -1162
rect 1490 -1193 1494 -1166
rect 1298 -1213 1325 -1209
rect 1310 -1231 1313 -1213
rect 1329 -1219 1332 -1205
rect 1422 -1208 1448 -1205
rect 1453 -1208 1457 -1197
rect 1476 -1208 1480 -1197
rect 1453 -1212 1480 -1208
rect 1467 -1231 1470 -1212
rect 1243 -1235 1470 -1231
rect 1484 -1240 1487 -1204
rect 1263 -1244 1487 -1240
rect 1098 -1252 1382 -1248
rect 1098 -1307 1104 -1252
rect 1115 -1259 1120 -1258
rect 1115 -1262 1328 -1259
rect 1115 -1263 1120 -1262
rect 1116 -1295 1119 -1263
rect 1163 -1280 1166 -1273
rect 1131 -1284 1225 -1280
rect 1138 -1290 1143 -1284
rect 1161 -1290 1166 -1284
rect 1199 -1290 1204 -1284
rect 1152 -1306 1156 -1296
rect 1175 -1306 1179 -1296
rect 1213 -1306 1217 -1296
rect 1098 -1311 1139 -1307
rect 1152 -1310 1200 -1306
rect 1213 -1310 1226 -1306
rect 1120 -1320 1162 -1316
rect 1175 -1327 1179 -1310
rect 1213 -1327 1217 -1310
rect 1156 -1332 1161 -1327
rect 1138 -1341 1142 -1332
rect 1199 -1341 1203 -1332
rect 1060 -1344 1199 -1341
rect 1223 -1362 1226 -1310
rect 1236 -1315 1241 -1262
rect 1259 -1306 1262 -1270
rect 1294 -1279 1297 -1273
rect 1271 -1283 1365 -1279
rect 1278 -1289 1283 -1283
rect 1301 -1289 1306 -1283
rect 1339 -1289 1344 -1283
rect 1292 -1305 1296 -1295
rect 1315 -1305 1319 -1295
rect 1353 -1305 1357 -1295
rect 1259 -1310 1279 -1306
rect 1292 -1309 1340 -1305
rect 1353 -1309 1364 -1305
rect 1236 -1319 1302 -1315
rect 1315 -1326 1319 -1309
rect 1353 -1326 1357 -1309
rect 1296 -1331 1301 -1326
rect 1278 -1340 1282 -1331
rect 1339 -1339 1343 -1331
rect 1278 -1341 1339 -1340
rect 1282 -1343 1339 -1341
rect 1361 -1350 1364 -1309
rect 1375 -1314 1382 -1252
rect 1397 -1305 1403 -1244
rect 1440 -1272 1603 -1269
rect 1436 -1278 1439 -1273
rect 1416 -1282 1510 -1278
rect 1598 -1279 1603 -1272
rect 1423 -1288 1428 -1282
rect 1446 -1288 1451 -1282
rect 1484 -1288 1489 -1282
rect 1584 -1283 1658 -1279
rect 1437 -1304 1441 -1294
rect 1460 -1304 1464 -1294
rect 1498 -1304 1502 -1294
rect 1584 -1291 1589 -1283
rect 1653 -1291 1658 -1283
rect 1602 -1297 1607 -1291
rect 1625 -1297 1630 -1291
rect 1397 -1309 1424 -1305
rect 1437 -1308 1485 -1304
rect 1498 -1308 1587 -1304
rect 1375 -1318 1447 -1314
rect 1460 -1325 1464 -1308
rect 1498 -1325 1502 -1308
rect 1644 -1309 1648 -1297
rect 1667 -1309 1671 -1297
rect 1644 -1313 1654 -1309
rect 1667 -1313 1681 -1309
rect 1644 -1314 1648 -1313
rect 1598 -1317 1648 -1314
rect 1598 -1320 1602 -1317
rect 1621 -1320 1625 -1317
rect 1644 -1320 1648 -1317
rect 1667 -1320 1671 -1313
rect 1441 -1330 1446 -1325
rect 1423 -1338 1427 -1330
rect 1484 -1338 1488 -1330
rect 1584 -1332 1588 -1325
rect 1607 -1332 1611 -1325
rect 1630 -1332 1634 -1325
rect 1653 -1332 1657 -1325
rect 1584 -1333 1657 -1332
rect 1504 -1336 1657 -1333
rect 1504 -1338 1509 -1336
rect 1484 -1339 1509 -1338
rect 1427 -1342 1509 -1339
rect 1513 -1345 1615 -1342
rect 1513 -1350 1517 -1345
rect 1361 -1354 1517 -1350
rect 1526 -1354 1637 -1350
rect 1526 -1362 1529 -1354
rect 1223 -1367 1529 -1362
rect 1676 -1403 1681 -1313
rect 878 -1418 1682 -1403
rect 1713 -1408 1722 -1118
rect 1894 -1267 1899 -1104
rect 2112 -1113 2161 -1109
rect 2112 -1138 2117 -1113
rect 1918 -1234 2064 -1230
rect 1918 -1340 1924 -1234
rect 2079 -1247 2082 -1167
rect 2112 -1193 2117 -1144
rect 2126 -1128 2148 -1123
rect 2126 -1138 2130 -1128
rect 2149 -1138 2153 -1128
rect 2126 -1193 2130 -1144
rect 2135 -1193 2140 -1144
rect 2149 -1193 2153 -1144
rect 2158 -1162 2161 -1113
rect 2173 -1121 2176 -1104
rect 2272 -1112 2316 -1108
rect 2166 -1126 2194 -1121
rect 2166 -1138 2171 -1126
rect 2189 -1138 2194 -1126
rect 2267 -1137 2272 -1113
rect 2161 -1166 2167 -1162
rect 2180 -1171 2184 -1144
rect 2158 -1175 2184 -1171
rect 2135 -1205 2140 -1197
rect 2158 -1205 2161 -1175
rect 2180 -1193 2184 -1175
rect 2203 -1162 2207 -1144
rect 2203 -1166 2216 -1162
rect 2203 -1193 2207 -1166
rect 2135 -1208 2161 -1205
rect 2267 -1192 2272 -1143
rect 2281 -1127 2308 -1122
rect 2281 -1137 2285 -1127
rect 2304 -1137 2308 -1127
rect 2281 -1192 2285 -1143
rect 2290 -1192 2295 -1143
rect 2304 -1192 2308 -1143
rect 2313 -1161 2316 -1112
rect 2332 -1120 2335 -1104
rect 2384 -1113 2389 -772
rect 2358 -1118 2389 -1113
rect 2321 -1125 2349 -1120
rect 2321 -1137 2326 -1125
rect 2344 -1137 2349 -1125
rect 2313 -1165 2322 -1161
rect 2335 -1170 2339 -1143
rect 2313 -1174 2339 -1170
rect 2166 -1208 2170 -1197
rect 2189 -1208 2193 -1197
rect 2290 -1204 2295 -1196
rect 2313 -1204 2316 -1174
rect 2335 -1192 2339 -1174
rect 2358 -1161 2362 -1143
rect 2358 -1165 2371 -1161
rect 2358 -1192 2362 -1165
rect 2166 -1212 2193 -1208
rect 2178 -1230 2181 -1212
rect 2197 -1218 2200 -1204
rect 2290 -1207 2316 -1204
rect 2321 -1207 2325 -1196
rect 2344 -1207 2348 -1196
rect 2321 -1211 2348 -1207
rect 2335 -1230 2338 -1211
rect 2111 -1234 2338 -1230
rect 2352 -1239 2355 -1203
rect 2131 -1243 2355 -1239
rect 1966 -1251 2250 -1247
rect 1966 -1306 1972 -1251
rect 1983 -1258 1988 -1257
rect 1983 -1261 2196 -1258
rect 1983 -1262 1988 -1261
rect 1984 -1294 1987 -1262
rect 2031 -1279 2034 -1272
rect 1999 -1283 2093 -1279
rect 2006 -1289 2011 -1283
rect 2029 -1289 2034 -1283
rect 2067 -1289 2072 -1283
rect 2020 -1305 2024 -1295
rect 2043 -1305 2047 -1295
rect 2081 -1305 2085 -1295
rect 1966 -1310 2007 -1306
rect 2020 -1309 2068 -1305
rect 2081 -1309 2094 -1305
rect 1988 -1319 2030 -1315
rect 2043 -1326 2047 -1309
rect 2081 -1326 2085 -1309
rect 2024 -1331 2029 -1326
rect 2006 -1340 2010 -1331
rect 2067 -1340 2071 -1331
rect 1928 -1343 2067 -1340
rect 2091 -1361 2094 -1309
rect 2104 -1314 2109 -1261
rect 2127 -1305 2130 -1269
rect 2162 -1278 2165 -1272
rect 2139 -1282 2233 -1278
rect 2146 -1288 2151 -1282
rect 2169 -1288 2174 -1282
rect 2207 -1288 2212 -1282
rect 2160 -1304 2164 -1294
rect 2183 -1304 2187 -1294
rect 2221 -1304 2225 -1294
rect 2127 -1309 2147 -1305
rect 2160 -1308 2208 -1304
rect 2221 -1308 2232 -1304
rect 2104 -1318 2170 -1314
rect 2183 -1325 2187 -1308
rect 2221 -1325 2225 -1308
rect 2164 -1330 2169 -1325
rect 2146 -1339 2150 -1330
rect 2207 -1338 2211 -1330
rect 2146 -1340 2207 -1339
rect 2150 -1342 2207 -1340
rect 2229 -1349 2232 -1308
rect 2243 -1313 2250 -1251
rect 2265 -1304 2271 -1243
rect 2308 -1271 2471 -1268
rect 2304 -1277 2307 -1272
rect 2284 -1281 2378 -1277
rect 2466 -1278 2471 -1271
rect 2291 -1287 2296 -1281
rect 2314 -1287 2319 -1281
rect 2352 -1287 2357 -1281
rect 2452 -1282 2526 -1278
rect 2305 -1303 2309 -1293
rect 2328 -1303 2332 -1293
rect 2366 -1303 2370 -1293
rect 2452 -1290 2457 -1282
rect 2521 -1290 2526 -1282
rect 2470 -1296 2475 -1290
rect 2493 -1296 2498 -1290
rect 2265 -1308 2292 -1304
rect 2305 -1307 2353 -1303
rect 2366 -1307 2455 -1303
rect 2243 -1317 2315 -1313
rect 2328 -1324 2332 -1307
rect 2366 -1324 2370 -1307
rect 2512 -1308 2516 -1296
rect 2535 -1308 2539 -1296
rect 2512 -1312 2522 -1308
rect 2535 -1312 2546 -1308
rect 2512 -1313 2516 -1312
rect 2466 -1316 2516 -1313
rect 2466 -1319 2470 -1316
rect 2489 -1319 2493 -1316
rect 2512 -1319 2516 -1316
rect 2535 -1319 2539 -1312
rect 2309 -1329 2314 -1324
rect 2291 -1337 2295 -1329
rect 2352 -1337 2356 -1329
rect 2452 -1331 2456 -1324
rect 2475 -1331 2479 -1324
rect 2498 -1331 2502 -1324
rect 2521 -1331 2525 -1324
rect 2452 -1332 2525 -1331
rect 2372 -1335 2525 -1332
rect 2372 -1337 2377 -1335
rect 2352 -1338 2377 -1337
rect 2295 -1341 2377 -1338
rect 2381 -1344 2483 -1341
rect 2381 -1349 2385 -1344
rect 2229 -1353 2385 -1349
rect 2394 -1353 2505 -1349
rect 2394 -1361 2397 -1353
rect 2091 -1366 2397 -1361
rect 2543 -1408 2546 -1312
rect 1713 -1418 2547 -1408
rect 1713 -1419 1902 -1418
rect -773 -1473 145 -1465
rect -765 -1475 145 -1473
rect 156 -1475 1049 -1465
rect 1060 -1475 1918 -1465
rect 1929 -1475 1932 -1465
<< m2contact >>
rect -771 -943 -760 -933
rect -460 -929 -455 -924
rect -687 -942 -676 -932
rect 330 -929 336 -924
rect 1311 -929 1318 -924
rect 2196 -928 2202 -923
rect 330 -949 336 -944
rect 1312 -948 1319 -943
rect -460 -957 -455 -952
rect 2195 -952 2204 -945
rect -494 -1170 -489 -1165
rect -678 -1275 -673 -1270
rect -508 -1237 -503 -1232
rect -424 -1131 -419 -1126
rect -305 -1116 -300 -1111
rect -416 -1170 -411 -1165
rect -466 -1237 -461 -1232
rect -376 -1226 -371 -1221
rect -446 -1246 -441 -1241
rect -376 -1264 -371 -1259
rect -542 -1275 -537 -1270
rect -589 -1302 -584 -1297
rect -589 -1323 -584 -1318
rect -505 -1348 -500 -1343
rect -446 -1272 -441 -1267
rect -411 -1275 -406 -1270
rect -427 -1348 -422 -1343
rect -365 -1346 -360 -1341
rect -269 -1275 -264 -1270
rect -282 -1345 -277 -1340
rect 307 -1168 312 -1163
rect 123 -1273 128 -1268
rect 293 -1235 298 -1230
rect 377 -1129 382 -1124
rect 496 -1114 501 -1109
rect 385 -1168 390 -1163
rect 335 -1235 340 -1230
rect 425 -1224 430 -1219
rect 355 -1244 360 -1239
rect 425 -1262 430 -1257
rect 259 -1273 264 -1268
rect 212 -1300 217 -1295
rect 212 -1321 217 -1316
rect 145 -1347 156 -1337
rect 296 -1346 301 -1341
rect 355 -1270 360 -1265
rect 390 -1273 395 -1268
rect 374 -1346 379 -1341
rect 436 -1344 441 -1339
rect 532 -1273 537 -1268
rect 519 -1343 524 -1338
rect 1210 -1168 1215 -1163
rect 1026 -1273 1031 -1268
rect 1196 -1235 1201 -1230
rect 1280 -1129 1285 -1124
rect 1399 -1114 1404 -1109
rect 1288 -1168 1293 -1163
rect 1238 -1235 1243 -1230
rect 1328 -1224 1333 -1219
rect 1258 -1244 1263 -1239
rect 1328 -1262 1333 -1257
rect 1162 -1273 1167 -1268
rect 1115 -1300 1120 -1295
rect 1115 -1321 1120 -1316
rect 1049 -1350 1060 -1340
rect 1199 -1346 1204 -1341
rect 1258 -1270 1263 -1265
rect 1293 -1273 1298 -1268
rect 1277 -1346 1282 -1341
rect 1339 -1344 1344 -1339
rect 1435 -1273 1440 -1268
rect 1422 -1343 1427 -1338
rect 2078 -1167 2083 -1162
rect 1894 -1272 1899 -1267
rect 2064 -1234 2069 -1229
rect 2148 -1128 2153 -1123
rect 2267 -1113 2272 -1108
rect 2156 -1167 2161 -1162
rect 2106 -1234 2111 -1229
rect 2196 -1223 2201 -1218
rect 2126 -1243 2131 -1238
rect 2196 -1261 2201 -1256
rect 2030 -1272 2035 -1267
rect 1983 -1299 1988 -1294
rect 1983 -1320 1988 -1315
rect 1918 -1349 1928 -1340
rect 2067 -1345 2072 -1340
rect 2126 -1269 2131 -1264
rect 2161 -1272 2166 -1267
rect 2145 -1345 2150 -1340
rect 2207 -1343 2212 -1338
rect 2303 -1272 2308 -1267
rect 2290 -1342 2295 -1337
rect 145 -1475 156 -1465
rect 1049 -1475 1060 -1465
rect 1918 -1475 1929 -1465
<< metal2 >>
rect -760 -942 -687 -934
rect -760 -943 -676 -942
rect -460 -952 -455 -929
rect 330 -944 335 -929
rect 1313 -943 1317 -929
rect 2197 -945 2201 -928
rect -344 -1115 -305 -1111
rect -344 -1118 -341 -1115
rect 457 -1113 496 -1109
rect 457 -1116 460 -1113
rect 1360 -1113 1399 -1109
rect 1360 -1116 1363 -1113
rect 2228 -1112 2267 -1108
rect 2228 -1115 2231 -1112
rect -423 -1122 -341 -1118
rect 378 -1120 460 -1116
rect 1281 -1120 1363 -1116
rect 2149 -1119 2231 -1115
rect -423 -1126 -420 -1122
rect 378 -1124 381 -1120
rect 1281 -1124 1284 -1120
rect 2149 -1123 2152 -1119
rect -489 -1169 -416 -1166
rect 312 -1167 385 -1164
rect 1215 -1167 1288 -1164
rect 2083 -1166 2156 -1163
rect -503 -1236 -466 -1233
rect -445 -1267 -442 -1246
rect -375 -1259 -372 -1226
rect 298 -1234 335 -1231
rect 356 -1265 359 -1244
rect 426 -1257 429 -1224
rect 1201 -1234 1238 -1231
rect 1259 -1265 1262 -1244
rect 1329 -1257 1332 -1224
rect 2069 -1233 2106 -1230
rect 2127 -1264 2130 -1243
rect 2197 -1256 2200 -1223
rect -673 -1274 -542 -1271
rect -537 -1274 -456 -1271
rect -459 -1277 -456 -1274
rect -432 -1274 -411 -1271
rect -432 -1277 -429 -1274
rect -406 -1274 -269 -1271
rect 128 -1272 259 -1269
rect 264 -1272 345 -1269
rect 342 -1275 345 -1272
rect 369 -1272 390 -1269
rect 369 -1275 372 -1272
rect 395 -1272 532 -1269
rect 1031 -1272 1162 -1269
rect 1167 -1272 1248 -1269
rect -459 -1280 -429 -1277
rect 342 -1278 372 -1275
rect 1245 -1275 1248 -1272
rect 1272 -1272 1293 -1269
rect 1272 -1275 1275 -1272
rect 1298 -1272 1435 -1269
rect 1899 -1271 2030 -1268
rect 2035 -1271 2116 -1268
rect 1245 -1278 1275 -1275
rect 2113 -1274 2116 -1271
rect 2140 -1271 2161 -1268
rect 2140 -1274 2143 -1271
rect 2166 -1271 2303 -1268
rect 2113 -1277 2143 -1274
rect -588 -1318 -585 -1302
rect 213 -1316 216 -1300
rect 1116 -1316 1119 -1300
rect 1984 -1315 1987 -1299
rect -500 -1347 -427 -1344
rect -360 -1345 -282 -1342
rect 301 -1345 374 -1342
rect 441 -1343 519 -1340
rect 145 -1465 155 -1347
rect 1204 -1345 1277 -1342
rect 1344 -1343 1422 -1340
rect 2072 -1344 2145 -1341
rect 2212 -1342 2290 -1339
rect 1049 -1465 1059 -1350
rect 1918 -1465 1928 -1349
<< labels >>
rlabel metal1 -322 -1106 -317 -1103 5 vdd
rlabel metal1 -309 -1237 -304 -1235 1 gnd
rlabel metal1 -32 -1314 -29 -1312 7 carry
rlabel polysilicon -399 -1168 -396 -1166 1 A3
rlabel polysilicon 402 -1167 406 -1163 1 A2
rlabel polysilicon 1305 -1167 1309 -1163 1 A1
rlabel polysilicon 2173 -1166 2177 -1162 1 A0
rlabel polysilicon -412 -858 -408 -854 1 B3
rlabel polysilicon 378 -858 382 -854 1 B2
rlabel polysilicon 1360 -858 1364 -854 1 B1
rlabel polysilicon 2244 -858 2248 -854 1 B0
rlabel metal1 2324 -771 2330 -769 1 M
rlabel metal1 -283 -1130 -276 -1126 1 Y3
rlabel metal1 519 -1128 526 -1124 1 Y2
rlabel metal1 1421 -1128 1428 -1124 1 Y1
rlabel metal1 2289 -1127 2296 -1123 1 Y0
<< end >>
