magic
tech scmos
timestamp 1700419032
<< nwell >>
rect 654 -5022 708 -5004
rect 715 -5022 746 -5004
rect 958 -5124 1012 -5106
rect 1019 -5124 1050 -5106
rect 1106 -5107 1137 -5089
rect 1196 -5120 1250 -5102
rect 1257 -5120 1288 -5102
rect 1327 -5120 1381 -5102
rect 1388 -5120 1419 -5102
rect 1483 -5120 1537 -5102
rect 1544 -5120 1575 -5102
rect 1105 -5175 1136 -5157
rect -591 -5339 -537 -5321
rect -525 -5339 -494 -5321
rect -483 -5339 -429 -5321
rect -417 -5339 -386 -5321
rect -371 -5339 -317 -5321
rect -305 -5339 -274 -5321
rect -259 -5339 -205 -5321
rect -193 -5339 -162 -5321
rect -148 -5339 -94 -5321
rect -82 -5339 -51 -5321
rect -36 -5339 18 -5321
rect 30 -5339 61 -5321
rect 76 -5339 130 -5321
rect 142 -5339 173 -5321
rect 188 -5339 242 -5321
rect 254 -5339 285 -5321
rect 560 -5332 614 -5314
rect 626 -5332 657 -5314
rect 668 -5332 722 -5314
rect 734 -5332 765 -5314
rect 780 -5332 834 -5314
rect 846 -5332 877 -5314
rect 892 -5332 946 -5314
rect 958 -5332 989 -5314
rect 1003 -5332 1057 -5314
rect 1069 -5332 1100 -5314
rect 1115 -5332 1169 -5314
rect 1181 -5332 1212 -5314
rect 1227 -5332 1281 -5314
rect 1293 -5332 1324 -5314
rect 1339 -5332 1393 -5314
rect 1405 -5332 1436 -5314
rect 1779 -5330 1833 -5312
rect 1845 -5330 1876 -5312
rect 1887 -5330 1941 -5312
rect 1953 -5330 1984 -5312
rect 1999 -5330 2053 -5312
rect 2065 -5330 2096 -5312
rect 2111 -5330 2165 -5312
rect 2177 -5330 2208 -5312
rect 2222 -5330 2276 -5312
rect 2288 -5330 2319 -5312
rect 2334 -5330 2388 -5312
rect 2400 -5330 2431 -5312
rect 2446 -5330 2500 -5312
rect 2512 -5330 2543 -5312
rect 2558 -5330 2612 -5312
rect 2624 -5330 2655 -5312
rect 2562 -5721 2685 -5703
rect -557 -5823 -503 -5805
rect -496 -5823 -465 -5805
rect -418 -5823 -364 -5805
rect -357 -5823 -326 -5805
rect -280 -5823 -226 -5805
rect -219 -5823 -188 -5805
rect -130 -5823 -76 -5805
rect -69 -5823 -38 -5805
rect 2087 -5870 2118 -5852
rect 2134 -5859 2188 -5841
rect 2213 -5859 2244 -5841
rect 2270 -5869 2301 -5851
rect 2335 -5859 2412 -5841
rect 2437 -5859 2468 -5841
rect 2498 -5869 2529 -5851
rect 2582 -5859 2682 -5841
rect 2707 -5859 2738 -5841
rect 2772 -5870 2803 -5852
rect 2862 -5859 2985 -5841
rect 3010 -5859 3041 -5841
rect 2076 -6002 2184 -5984
rect 2210 -6007 2241 -5989
rect 2075 -6147 2183 -6129
rect 2209 -6152 2240 -6134
rect -1589 -6180 -1481 -6162
rect -799 -6180 -691 -6162
rect 183 -6180 291 -6162
rect 1067 -6180 1175 -6162
rect 2339 -6234 2439 -6216
rect 2464 -6234 2495 -6216
rect 2075 -6309 2183 -6291
rect 2209 -6314 2240 -6296
rect 2076 -6463 2184 -6445
rect 2210 -6468 2241 -6450
rect -1576 -6491 -1468 -6473
rect -1421 -6490 -1313 -6472
rect -775 -6489 -667 -6471
rect -620 -6488 -512 -6470
rect 128 -6489 236 -6471
rect 283 -6488 391 -6470
rect 996 -6488 1104 -6470
rect 1151 -6487 1259 -6469
rect -1682 -6642 -1628 -6624
rect -1621 -6642 -1590 -6624
rect -1542 -6641 -1488 -6623
rect -1481 -6641 -1450 -6623
rect -1397 -6640 -1343 -6622
rect -1336 -6640 -1305 -6622
rect -1236 -6643 -1136 -6625
rect -881 -6640 -827 -6622
rect -820 -6640 -789 -6622
rect -741 -6639 -687 -6621
rect -680 -6639 -649 -6621
rect -596 -6638 -542 -6620
rect -535 -6638 -504 -6620
rect -435 -6641 -335 -6623
rect 22 -6640 76 -6622
rect 83 -6640 114 -6622
rect 162 -6639 216 -6621
rect 223 -6639 254 -6621
rect 307 -6638 361 -6620
rect 368 -6638 399 -6620
rect 468 -6641 568 -6623
rect 890 -6639 944 -6621
rect 951 -6639 982 -6621
rect 1030 -6638 1084 -6620
rect 1091 -6638 1122 -6620
rect 1175 -6637 1229 -6619
rect 1236 -6637 1267 -6619
rect 1336 -6640 1436 -6622
rect 2081 -6678 2112 -6660
rect 2128 -6667 2182 -6649
rect 2207 -6667 2238 -6649
rect 2272 -6677 2303 -6659
rect 2337 -6667 2414 -6649
rect 2439 -6667 2470 -6649
rect 2499 -6677 2530 -6659
rect 2583 -6667 2683 -6649
rect 2708 -6667 2739 -6649
rect 2770 -6677 2801 -6659
rect 2860 -6666 2983 -6648
rect 3008 -6666 3039 -6648
rect 3092 -6660 3215 -6642
<< ntransistor >>
rect 669 -5052 672 -5047
rect 692 -5052 695 -5047
rect 730 -5052 733 -5047
rect 1121 -5127 1124 -5122
rect 973 -5154 976 -5149
rect 996 -5154 999 -5149
rect 1034 -5154 1037 -5149
rect 1211 -5150 1214 -5145
rect 1234 -5150 1237 -5145
rect 1272 -5150 1275 -5145
rect 1342 -5150 1345 -5145
rect 1365 -5150 1368 -5145
rect 1403 -5150 1406 -5145
rect 1498 -5150 1501 -5145
rect 1521 -5150 1524 -5145
rect 1559 -5150 1562 -5145
rect 1120 -5195 1123 -5190
rect 575 -5362 578 -5357
rect 598 -5362 601 -5357
rect 641 -5362 644 -5357
rect 683 -5362 686 -5357
rect 706 -5362 709 -5357
rect 749 -5362 752 -5357
rect 795 -5362 798 -5357
rect 818 -5362 821 -5357
rect 861 -5362 864 -5357
rect 907 -5362 910 -5357
rect 930 -5362 933 -5357
rect 973 -5362 976 -5357
rect 1018 -5362 1021 -5357
rect 1041 -5362 1044 -5357
rect 1084 -5362 1087 -5357
rect 1130 -5362 1133 -5357
rect 1153 -5362 1156 -5357
rect 1196 -5362 1199 -5357
rect 1242 -5362 1245 -5357
rect 1265 -5362 1268 -5357
rect 1308 -5362 1311 -5357
rect 1354 -5362 1357 -5357
rect 1377 -5362 1380 -5357
rect 1420 -5362 1423 -5357
rect 1794 -5360 1797 -5355
rect 1817 -5360 1820 -5355
rect 1860 -5360 1863 -5355
rect 1902 -5360 1905 -5355
rect 1925 -5360 1928 -5355
rect 1968 -5360 1971 -5355
rect 2014 -5360 2017 -5355
rect 2037 -5360 2040 -5355
rect 2080 -5360 2083 -5355
rect 2126 -5360 2129 -5355
rect 2149 -5360 2152 -5355
rect 2192 -5360 2195 -5355
rect 2237 -5360 2240 -5355
rect 2260 -5360 2263 -5355
rect 2303 -5360 2306 -5355
rect 2349 -5360 2352 -5355
rect 2372 -5360 2375 -5355
rect 2415 -5360 2418 -5355
rect 2461 -5360 2464 -5355
rect 2484 -5360 2487 -5355
rect 2527 -5360 2530 -5355
rect 2573 -5360 2576 -5355
rect 2596 -5360 2599 -5355
rect 2639 -5360 2642 -5355
rect -576 -5369 -573 -5364
rect -553 -5369 -550 -5364
rect -510 -5369 -507 -5364
rect -468 -5369 -465 -5364
rect -445 -5369 -442 -5364
rect -402 -5369 -399 -5364
rect -356 -5369 -353 -5364
rect -333 -5369 -330 -5364
rect -290 -5369 -287 -5364
rect -244 -5369 -241 -5364
rect -221 -5369 -218 -5364
rect -178 -5369 -175 -5364
rect -133 -5369 -130 -5364
rect -110 -5369 -107 -5364
rect -67 -5369 -64 -5364
rect -21 -5369 -18 -5364
rect 2 -5369 5 -5364
rect 45 -5369 48 -5364
rect 91 -5369 94 -5364
rect 114 -5369 117 -5364
rect 157 -5369 160 -5364
rect 203 -5369 206 -5364
rect 226 -5369 229 -5364
rect 269 -5369 272 -5364
rect 2577 -5743 2580 -5738
rect 2600 -5743 2603 -5738
rect 2623 -5743 2626 -5738
rect 2646 -5743 2649 -5738
rect 2669 -5743 2672 -5738
rect -542 -5853 -539 -5848
rect -519 -5853 -516 -5848
rect -481 -5853 -478 -5848
rect -403 -5853 -400 -5848
rect -380 -5853 -377 -5848
rect -342 -5853 -339 -5848
rect -265 -5853 -262 -5848
rect -242 -5853 -239 -5848
rect -204 -5853 -201 -5848
rect -115 -5853 -112 -5848
rect -92 -5853 -89 -5848
rect -54 -5853 -51 -5848
rect 2102 -5890 2105 -5885
rect 2149 -5889 2152 -5884
rect 2172 -5889 2175 -5884
rect 2228 -5889 2231 -5884
rect 2285 -5889 2288 -5884
rect 2350 -5889 2353 -5884
rect 2373 -5889 2376 -5884
rect 2396 -5889 2399 -5884
rect 2452 -5889 2455 -5884
rect 2513 -5889 2516 -5884
rect 2597 -5889 2600 -5884
rect 2620 -5889 2623 -5884
rect 2643 -5889 2646 -5884
rect 2666 -5889 2669 -5884
rect 2722 -5889 2725 -5884
rect 2787 -5890 2790 -5885
rect 2877 -5889 2880 -5884
rect 2900 -5889 2903 -5884
rect 2923 -5889 2926 -5884
rect 2946 -5889 2949 -5884
rect 2969 -5889 2972 -5884
rect 3025 -5889 3028 -5884
rect 2091 -6049 2094 -6045
rect 2114 -6049 2117 -6045
rect 2145 -6049 2148 -6045
rect 2168 -6049 2171 -6045
rect 2225 -6027 2228 -6022
rect -1574 -6227 -1571 -6223
rect -1551 -6227 -1548 -6223
rect -1520 -6227 -1517 -6223
rect -1497 -6227 -1494 -6223
rect -784 -6227 -781 -6223
rect -761 -6227 -758 -6223
rect -730 -6227 -727 -6223
rect -707 -6227 -704 -6223
rect 198 -6227 201 -6223
rect 221 -6227 224 -6223
rect 252 -6227 255 -6223
rect 275 -6227 278 -6223
rect 1082 -6227 1085 -6223
rect 1105 -6227 1108 -6223
rect 1136 -6227 1139 -6223
rect 1159 -6227 1162 -6223
rect 2090 -6194 2093 -6190
rect 2113 -6194 2116 -6190
rect 2144 -6194 2147 -6190
rect 2167 -6194 2170 -6190
rect 2224 -6172 2227 -6167
rect 2354 -6264 2357 -6259
rect 2377 -6264 2380 -6259
rect 2400 -6264 2403 -6259
rect 2423 -6264 2426 -6259
rect 2479 -6264 2482 -6259
rect 2090 -6356 2093 -6352
rect 2113 -6356 2116 -6352
rect 2144 -6356 2147 -6352
rect 2167 -6356 2170 -6352
rect 2224 -6334 2227 -6329
rect -1561 -6538 -1558 -6534
rect -1538 -6538 -1535 -6534
rect -1507 -6538 -1504 -6534
rect -1484 -6538 -1481 -6534
rect -1406 -6537 -1403 -6533
rect -1383 -6537 -1380 -6533
rect -1352 -6537 -1349 -6533
rect -1329 -6537 -1326 -6533
rect -760 -6536 -757 -6532
rect -737 -6536 -734 -6532
rect -706 -6536 -703 -6532
rect -683 -6536 -680 -6532
rect -605 -6535 -602 -6531
rect -582 -6535 -579 -6531
rect -551 -6535 -548 -6531
rect -528 -6535 -525 -6531
rect 143 -6536 146 -6532
rect 166 -6536 169 -6532
rect 197 -6536 200 -6532
rect 220 -6536 223 -6532
rect 298 -6535 301 -6531
rect 321 -6535 324 -6531
rect 352 -6535 355 -6531
rect 375 -6535 378 -6531
rect 1011 -6535 1014 -6531
rect 1034 -6535 1037 -6531
rect 1065 -6535 1068 -6531
rect 1088 -6535 1091 -6531
rect 1166 -6534 1169 -6530
rect 1189 -6534 1192 -6530
rect 1220 -6534 1223 -6530
rect 1243 -6534 1246 -6530
rect 2091 -6510 2094 -6506
rect 2114 -6510 2117 -6506
rect 2145 -6510 2148 -6506
rect 2168 -6510 2171 -6506
rect 2225 -6488 2228 -6483
rect -1221 -6665 -1218 -6660
rect -1198 -6665 -1195 -6660
rect -1175 -6665 -1172 -6660
rect -1152 -6665 -1149 -6660
rect -420 -6663 -417 -6658
rect -397 -6663 -394 -6658
rect -374 -6663 -371 -6658
rect -351 -6663 -348 -6658
rect -1667 -6672 -1664 -6667
rect -1644 -6672 -1641 -6667
rect -1606 -6672 -1603 -6667
rect -1527 -6671 -1524 -6666
rect -1504 -6671 -1501 -6666
rect -1466 -6671 -1463 -6666
rect -1382 -6670 -1379 -6665
rect -1359 -6670 -1356 -6665
rect -1321 -6670 -1318 -6665
rect -866 -6670 -863 -6665
rect -843 -6670 -840 -6665
rect -805 -6670 -802 -6665
rect -726 -6669 -723 -6664
rect -703 -6669 -700 -6664
rect -665 -6669 -662 -6664
rect -581 -6668 -578 -6663
rect -558 -6668 -555 -6663
rect -520 -6668 -517 -6663
rect 483 -6663 486 -6658
rect 506 -6663 509 -6658
rect 529 -6663 532 -6658
rect 552 -6663 555 -6658
rect 37 -6670 40 -6665
rect 60 -6670 63 -6665
rect 98 -6670 101 -6665
rect 177 -6669 180 -6664
rect 200 -6669 203 -6664
rect 238 -6669 241 -6664
rect 322 -6668 325 -6663
rect 345 -6668 348 -6663
rect 383 -6668 386 -6663
rect 1351 -6662 1354 -6657
rect 1374 -6662 1377 -6657
rect 1397 -6662 1400 -6657
rect 1420 -6662 1423 -6657
rect 905 -6669 908 -6664
rect 928 -6669 931 -6664
rect 966 -6669 969 -6664
rect 1045 -6668 1048 -6663
rect 1068 -6668 1071 -6663
rect 1106 -6668 1109 -6663
rect 1190 -6667 1193 -6662
rect 1213 -6667 1216 -6662
rect 1251 -6667 1254 -6662
rect 3107 -6682 3110 -6677
rect 3130 -6682 3133 -6677
rect 3153 -6682 3156 -6677
rect 3176 -6682 3179 -6677
rect 3199 -6682 3202 -6677
rect 2096 -6698 2099 -6693
rect 2143 -6697 2146 -6692
rect 2166 -6697 2169 -6692
rect 2222 -6697 2225 -6692
rect 2287 -6697 2290 -6692
rect 2352 -6697 2355 -6692
rect 2375 -6697 2378 -6692
rect 2398 -6697 2401 -6692
rect 2454 -6697 2457 -6692
rect 2514 -6697 2517 -6692
rect 2598 -6697 2601 -6692
rect 2621 -6697 2624 -6692
rect 2644 -6697 2647 -6692
rect 2667 -6697 2670 -6692
rect 2723 -6697 2726 -6692
rect 2785 -6697 2788 -6692
rect 2875 -6696 2878 -6691
rect 2898 -6696 2901 -6691
rect 2921 -6696 2924 -6691
rect 2944 -6696 2947 -6691
rect 2967 -6696 2970 -6691
rect 3023 -6696 3026 -6691
<< ptransistor >>
rect 669 -5016 672 -5010
rect 692 -5016 695 -5010
rect 730 -5016 733 -5010
rect 1121 -5101 1124 -5095
rect 973 -5118 976 -5112
rect 996 -5118 999 -5112
rect 1034 -5118 1037 -5112
rect 1211 -5114 1214 -5108
rect 1234 -5114 1237 -5108
rect 1272 -5114 1275 -5108
rect 1342 -5114 1345 -5108
rect 1365 -5114 1368 -5108
rect 1403 -5114 1406 -5108
rect 1498 -5114 1501 -5108
rect 1521 -5114 1524 -5108
rect 1559 -5114 1562 -5108
rect 1120 -5169 1123 -5163
rect 575 -5326 578 -5320
rect 598 -5326 601 -5320
rect 641 -5326 644 -5320
rect 683 -5326 686 -5320
rect 706 -5326 709 -5320
rect 749 -5326 752 -5320
rect 795 -5326 798 -5320
rect 818 -5326 821 -5320
rect 861 -5326 864 -5320
rect 907 -5326 910 -5320
rect 930 -5326 933 -5320
rect 973 -5326 976 -5320
rect 1018 -5326 1021 -5320
rect 1041 -5326 1044 -5320
rect 1084 -5326 1087 -5320
rect 1130 -5326 1133 -5320
rect 1153 -5326 1156 -5320
rect 1196 -5326 1199 -5320
rect 1242 -5326 1245 -5320
rect 1265 -5326 1268 -5320
rect 1308 -5326 1311 -5320
rect 1354 -5326 1357 -5320
rect 1377 -5326 1380 -5320
rect 1420 -5326 1423 -5320
rect 1794 -5324 1797 -5318
rect 1817 -5324 1820 -5318
rect 1860 -5324 1863 -5318
rect 1902 -5324 1905 -5318
rect 1925 -5324 1928 -5318
rect 1968 -5324 1971 -5318
rect 2014 -5324 2017 -5318
rect 2037 -5324 2040 -5318
rect 2080 -5324 2083 -5318
rect 2126 -5324 2129 -5318
rect 2149 -5324 2152 -5318
rect 2192 -5324 2195 -5318
rect 2237 -5324 2240 -5318
rect 2260 -5324 2263 -5318
rect 2303 -5324 2306 -5318
rect 2349 -5324 2352 -5318
rect 2372 -5324 2375 -5318
rect 2415 -5324 2418 -5318
rect 2461 -5324 2464 -5318
rect 2484 -5324 2487 -5318
rect 2527 -5324 2530 -5318
rect 2573 -5324 2576 -5318
rect 2596 -5324 2599 -5318
rect 2639 -5324 2642 -5318
rect -576 -5333 -573 -5327
rect -553 -5333 -550 -5327
rect -510 -5333 -507 -5327
rect -468 -5333 -465 -5327
rect -445 -5333 -442 -5327
rect -402 -5333 -399 -5327
rect -356 -5333 -353 -5327
rect -333 -5333 -330 -5327
rect -290 -5333 -287 -5327
rect -244 -5333 -241 -5327
rect -221 -5333 -218 -5327
rect -178 -5333 -175 -5327
rect -133 -5333 -130 -5327
rect -110 -5333 -107 -5327
rect -67 -5333 -64 -5327
rect -21 -5333 -18 -5327
rect 2 -5333 5 -5327
rect 45 -5333 48 -5327
rect 91 -5333 94 -5327
rect 114 -5333 117 -5327
rect 157 -5333 160 -5327
rect 203 -5333 206 -5327
rect 226 -5333 229 -5327
rect 269 -5333 272 -5327
rect 2577 -5715 2580 -5709
rect 2600 -5715 2603 -5709
rect 2623 -5715 2626 -5709
rect 2646 -5715 2649 -5709
rect 2669 -5715 2672 -5709
rect -542 -5817 -539 -5811
rect -519 -5817 -516 -5811
rect -481 -5817 -478 -5811
rect -403 -5817 -400 -5811
rect -380 -5817 -377 -5811
rect -342 -5817 -339 -5811
rect -265 -5817 -262 -5811
rect -242 -5817 -239 -5811
rect -204 -5817 -201 -5811
rect -115 -5817 -112 -5811
rect -92 -5817 -89 -5811
rect -54 -5817 -51 -5811
rect 2149 -5853 2152 -5847
rect 2172 -5853 2175 -5847
rect 2228 -5853 2231 -5847
rect 2350 -5853 2353 -5847
rect 2373 -5853 2376 -5847
rect 2396 -5853 2399 -5847
rect 2452 -5853 2455 -5847
rect 2597 -5853 2600 -5847
rect 2620 -5853 2623 -5847
rect 2643 -5853 2646 -5847
rect 2666 -5853 2669 -5847
rect 2722 -5853 2725 -5847
rect 2877 -5853 2880 -5847
rect 2900 -5853 2903 -5847
rect 2923 -5853 2926 -5847
rect 2946 -5853 2949 -5847
rect 2969 -5853 2972 -5847
rect 3025 -5853 3028 -5847
rect 2102 -5864 2105 -5858
rect 2285 -5863 2288 -5857
rect 2513 -5863 2516 -5857
rect 2787 -5864 2790 -5858
rect 2091 -5996 2094 -5990
rect 2114 -5996 2117 -5990
rect 2145 -5996 2148 -5990
rect 2168 -5996 2171 -5990
rect 2225 -6001 2228 -5995
rect -1574 -6174 -1571 -6168
rect -1551 -6174 -1548 -6168
rect -1520 -6174 -1517 -6168
rect -1497 -6174 -1494 -6168
rect -784 -6174 -781 -6168
rect -761 -6174 -758 -6168
rect -730 -6174 -727 -6168
rect -707 -6174 -704 -6168
rect 198 -6174 201 -6168
rect 221 -6174 224 -6168
rect 252 -6174 255 -6168
rect 275 -6174 278 -6168
rect 1082 -6174 1085 -6168
rect 1105 -6174 1108 -6168
rect 1136 -6174 1139 -6168
rect 1159 -6174 1162 -6168
rect 2090 -6141 2093 -6135
rect 2113 -6141 2116 -6135
rect 2144 -6141 2147 -6135
rect 2167 -6141 2170 -6135
rect 2224 -6146 2227 -6140
rect 2354 -6228 2357 -6222
rect 2377 -6228 2380 -6222
rect 2400 -6228 2403 -6222
rect 2423 -6228 2426 -6222
rect 2479 -6228 2482 -6222
rect 2090 -6303 2093 -6297
rect 2113 -6303 2116 -6297
rect 2144 -6303 2147 -6297
rect 2167 -6303 2170 -6297
rect 2224 -6308 2227 -6302
rect -1561 -6485 -1558 -6479
rect -1538 -6485 -1535 -6479
rect -1507 -6485 -1504 -6479
rect -1484 -6485 -1481 -6479
rect -1406 -6484 -1403 -6478
rect -1383 -6484 -1380 -6478
rect -1352 -6484 -1349 -6478
rect -1329 -6484 -1326 -6478
rect -760 -6483 -757 -6477
rect -737 -6483 -734 -6477
rect -706 -6483 -703 -6477
rect -683 -6483 -680 -6477
rect -605 -6482 -602 -6476
rect -582 -6482 -579 -6476
rect -551 -6482 -548 -6476
rect -528 -6482 -525 -6476
rect 143 -6483 146 -6477
rect 166 -6483 169 -6477
rect 197 -6483 200 -6477
rect 220 -6483 223 -6477
rect 298 -6482 301 -6476
rect 321 -6482 324 -6476
rect 352 -6482 355 -6476
rect 375 -6482 378 -6476
rect 1011 -6482 1014 -6476
rect 1034 -6482 1037 -6476
rect 1065 -6482 1068 -6476
rect 1088 -6482 1091 -6476
rect 1166 -6481 1169 -6475
rect 1189 -6481 1192 -6475
rect 1220 -6481 1223 -6475
rect 1243 -6481 1246 -6475
rect 2091 -6457 2094 -6451
rect 2114 -6457 2117 -6451
rect 2145 -6457 2148 -6451
rect 2168 -6457 2171 -6451
rect 2225 -6462 2228 -6456
rect -1667 -6636 -1664 -6630
rect -1644 -6636 -1641 -6630
rect -1606 -6636 -1603 -6630
rect -1527 -6635 -1524 -6629
rect -1504 -6635 -1501 -6629
rect -1466 -6635 -1463 -6629
rect -1382 -6634 -1379 -6628
rect -1359 -6634 -1356 -6628
rect -1321 -6634 -1318 -6628
rect -1221 -6637 -1218 -6631
rect -1198 -6637 -1195 -6631
rect -1175 -6637 -1172 -6631
rect -1152 -6637 -1149 -6631
rect -866 -6634 -863 -6628
rect -843 -6634 -840 -6628
rect -805 -6634 -802 -6628
rect -726 -6633 -723 -6627
rect -703 -6633 -700 -6627
rect -665 -6633 -662 -6627
rect -581 -6632 -578 -6626
rect -558 -6632 -555 -6626
rect -520 -6632 -517 -6626
rect -420 -6635 -417 -6629
rect -397 -6635 -394 -6629
rect -374 -6635 -371 -6629
rect -351 -6635 -348 -6629
rect 37 -6634 40 -6628
rect 60 -6634 63 -6628
rect 98 -6634 101 -6628
rect 177 -6633 180 -6627
rect 200 -6633 203 -6627
rect 238 -6633 241 -6627
rect 322 -6632 325 -6626
rect 345 -6632 348 -6626
rect 383 -6632 386 -6626
rect 483 -6635 486 -6629
rect 506 -6635 509 -6629
rect 529 -6635 532 -6629
rect 552 -6635 555 -6629
rect 905 -6633 908 -6627
rect 928 -6633 931 -6627
rect 966 -6633 969 -6627
rect 1045 -6632 1048 -6626
rect 1068 -6632 1071 -6626
rect 1106 -6632 1109 -6626
rect 1190 -6631 1193 -6625
rect 1213 -6631 1216 -6625
rect 1251 -6631 1254 -6625
rect 1351 -6634 1354 -6628
rect 1374 -6634 1377 -6628
rect 1397 -6634 1400 -6628
rect 1420 -6634 1423 -6628
rect 3107 -6654 3110 -6648
rect 3130 -6654 3133 -6648
rect 3153 -6654 3156 -6648
rect 3176 -6654 3179 -6648
rect 3199 -6654 3202 -6648
rect 2143 -6661 2146 -6655
rect 2166 -6661 2169 -6655
rect 2222 -6661 2225 -6655
rect 2352 -6661 2355 -6655
rect 2375 -6661 2378 -6655
rect 2398 -6661 2401 -6655
rect 2454 -6661 2457 -6655
rect 2598 -6661 2601 -6655
rect 2621 -6661 2624 -6655
rect 2644 -6661 2647 -6655
rect 2667 -6661 2670 -6655
rect 2723 -6661 2726 -6655
rect 2875 -6660 2878 -6654
rect 2898 -6660 2901 -6654
rect 2921 -6660 2924 -6654
rect 2944 -6660 2947 -6654
rect 2967 -6660 2970 -6654
rect 3023 -6660 3026 -6654
rect 2096 -6672 2099 -6666
rect 2287 -6671 2290 -6665
rect 2514 -6671 2517 -6665
rect 2785 -6671 2788 -6665
<< ndiffusion >>
rect 665 -5052 669 -5047
rect 672 -5052 675 -5047
rect 688 -5052 692 -5047
rect 695 -5052 698 -5047
rect 726 -5052 730 -5047
rect 733 -5052 736 -5047
rect 1117 -5127 1121 -5122
rect 1124 -5127 1127 -5122
rect 969 -5154 973 -5149
rect 976 -5154 979 -5149
rect 992 -5154 996 -5149
rect 999 -5154 1002 -5149
rect 1030 -5154 1034 -5149
rect 1037 -5154 1040 -5149
rect 1207 -5150 1211 -5145
rect 1214 -5150 1217 -5145
rect 1230 -5150 1234 -5145
rect 1237 -5150 1240 -5145
rect 1268 -5150 1272 -5145
rect 1275 -5150 1278 -5145
rect 1338 -5150 1342 -5145
rect 1345 -5150 1348 -5145
rect 1361 -5150 1365 -5145
rect 1368 -5150 1371 -5145
rect 1399 -5150 1403 -5145
rect 1406 -5150 1409 -5145
rect 1494 -5150 1498 -5145
rect 1501 -5150 1504 -5145
rect 1517 -5150 1521 -5145
rect 1524 -5150 1527 -5145
rect 1555 -5150 1559 -5145
rect 1562 -5150 1565 -5145
rect 1116 -5195 1120 -5190
rect 1123 -5195 1126 -5190
rect 571 -5362 575 -5357
rect 578 -5362 581 -5357
rect 594 -5362 598 -5357
rect 601 -5362 604 -5357
rect 637 -5362 641 -5357
rect 644 -5362 647 -5357
rect 679 -5362 683 -5357
rect 686 -5362 689 -5357
rect 702 -5362 706 -5357
rect 709 -5362 712 -5357
rect 745 -5362 749 -5357
rect 752 -5362 755 -5357
rect 791 -5362 795 -5357
rect 798 -5362 801 -5357
rect 814 -5362 818 -5357
rect 821 -5362 824 -5357
rect 857 -5362 861 -5357
rect 864 -5362 867 -5357
rect 903 -5362 907 -5357
rect 910 -5362 913 -5357
rect 926 -5362 930 -5357
rect 933 -5362 936 -5357
rect 969 -5362 973 -5357
rect 976 -5362 979 -5357
rect 1014 -5362 1018 -5357
rect 1021 -5362 1024 -5357
rect 1037 -5362 1041 -5357
rect 1044 -5362 1047 -5357
rect 1080 -5362 1084 -5357
rect 1087 -5362 1090 -5357
rect 1126 -5362 1130 -5357
rect 1133 -5362 1136 -5357
rect 1149 -5362 1153 -5357
rect 1156 -5362 1159 -5357
rect 1192 -5362 1196 -5357
rect 1199 -5362 1202 -5357
rect 1238 -5362 1242 -5357
rect 1245 -5362 1248 -5357
rect 1261 -5362 1265 -5357
rect 1268 -5362 1271 -5357
rect 1304 -5362 1308 -5357
rect 1311 -5362 1314 -5357
rect 1350 -5362 1354 -5357
rect 1357 -5362 1360 -5357
rect 1373 -5362 1377 -5357
rect 1380 -5362 1383 -5357
rect 1416 -5362 1420 -5357
rect 1423 -5362 1426 -5357
rect 1790 -5360 1794 -5355
rect 1797 -5360 1800 -5355
rect 1813 -5360 1817 -5355
rect 1820 -5360 1823 -5355
rect 1856 -5360 1860 -5355
rect 1863 -5360 1866 -5355
rect 1898 -5360 1902 -5355
rect 1905 -5360 1908 -5355
rect 1921 -5360 1925 -5355
rect 1928 -5360 1931 -5355
rect 1964 -5360 1968 -5355
rect 1971 -5360 1974 -5355
rect 2010 -5360 2014 -5355
rect 2017 -5360 2020 -5355
rect 2033 -5360 2037 -5355
rect 2040 -5360 2043 -5355
rect 2076 -5360 2080 -5355
rect 2083 -5360 2086 -5355
rect 2122 -5360 2126 -5355
rect 2129 -5360 2132 -5355
rect 2145 -5360 2149 -5355
rect 2152 -5360 2155 -5355
rect 2188 -5360 2192 -5355
rect 2195 -5360 2198 -5355
rect 2233 -5360 2237 -5355
rect 2240 -5360 2243 -5355
rect 2256 -5360 2260 -5355
rect 2263 -5360 2266 -5355
rect 2299 -5360 2303 -5355
rect 2306 -5360 2309 -5355
rect 2345 -5360 2349 -5355
rect 2352 -5360 2355 -5355
rect 2368 -5360 2372 -5355
rect 2375 -5360 2378 -5355
rect 2411 -5360 2415 -5355
rect 2418 -5360 2421 -5355
rect 2457 -5360 2461 -5355
rect 2464 -5360 2467 -5355
rect 2480 -5360 2484 -5355
rect 2487 -5360 2490 -5355
rect 2523 -5360 2527 -5355
rect 2530 -5360 2533 -5355
rect 2569 -5360 2573 -5355
rect 2576 -5360 2579 -5355
rect 2592 -5360 2596 -5355
rect 2599 -5360 2602 -5355
rect 2635 -5360 2639 -5355
rect 2642 -5360 2645 -5355
rect -580 -5369 -576 -5364
rect -573 -5369 -570 -5364
rect -557 -5369 -553 -5364
rect -550 -5369 -547 -5364
rect -514 -5369 -510 -5364
rect -507 -5369 -504 -5364
rect -472 -5369 -468 -5364
rect -465 -5369 -462 -5364
rect -449 -5369 -445 -5364
rect -442 -5369 -439 -5364
rect -406 -5369 -402 -5364
rect -399 -5369 -396 -5364
rect -360 -5369 -356 -5364
rect -353 -5369 -350 -5364
rect -337 -5369 -333 -5364
rect -330 -5369 -327 -5364
rect -294 -5369 -290 -5364
rect -287 -5369 -284 -5364
rect -248 -5369 -244 -5364
rect -241 -5369 -238 -5364
rect -225 -5369 -221 -5364
rect -218 -5369 -215 -5364
rect -182 -5369 -178 -5364
rect -175 -5369 -172 -5364
rect -137 -5369 -133 -5364
rect -130 -5369 -127 -5364
rect -114 -5369 -110 -5364
rect -107 -5369 -104 -5364
rect -71 -5369 -67 -5364
rect -64 -5369 -61 -5364
rect -25 -5369 -21 -5364
rect -18 -5369 -15 -5364
rect -2 -5369 2 -5364
rect 5 -5369 8 -5364
rect 41 -5369 45 -5364
rect 48 -5369 51 -5364
rect 87 -5369 91 -5364
rect 94 -5369 97 -5364
rect 110 -5369 114 -5364
rect 117 -5369 120 -5364
rect 153 -5369 157 -5364
rect 160 -5369 163 -5364
rect 199 -5369 203 -5364
rect 206 -5369 209 -5364
rect 222 -5369 226 -5364
rect 229 -5369 232 -5364
rect 265 -5369 269 -5364
rect 272 -5369 275 -5364
rect 2573 -5743 2577 -5738
rect 2580 -5743 2583 -5738
rect 2596 -5743 2600 -5738
rect 2603 -5743 2606 -5738
rect 2619 -5743 2623 -5738
rect 2626 -5743 2629 -5738
rect 2642 -5743 2646 -5738
rect 2649 -5743 2652 -5738
rect 2665 -5743 2669 -5738
rect 2672 -5743 2675 -5738
rect -546 -5853 -542 -5848
rect -539 -5853 -536 -5848
rect -523 -5853 -519 -5848
rect -516 -5853 -513 -5848
rect -485 -5853 -481 -5848
rect -478 -5853 -475 -5848
rect -407 -5853 -403 -5848
rect -400 -5853 -397 -5848
rect -384 -5853 -380 -5848
rect -377 -5853 -374 -5848
rect -346 -5853 -342 -5848
rect -339 -5853 -336 -5848
rect -269 -5853 -265 -5848
rect -262 -5853 -259 -5848
rect -246 -5853 -242 -5848
rect -239 -5853 -236 -5848
rect -208 -5853 -204 -5848
rect -201 -5853 -198 -5848
rect -119 -5853 -115 -5848
rect -112 -5853 -109 -5848
rect -96 -5853 -92 -5848
rect -89 -5853 -86 -5848
rect -58 -5853 -54 -5848
rect -51 -5853 -48 -5848
rect 2098 -5890 2102 -5885
rect 2105 -5890 2108 -5885
rect 2145 -5889 2149 -5884
rect 2152 -5889 2155 -5884
rect 2168 -5889 2172 -5884
rect 2175 -5889 2178 -5884
rect 2224 -5889 2228 -5884
rect 2231 -5889 2234 -5884
rect 2281 -5889 2285 -5884
rect 2288 -5889 2291 -5884
rect 2346 -5889 2350 -5884
rect 2353 -5889 2356 -5884
rect 2369 -5889 2373 -5884
rect 2376 -5889 2379 -5884
rect 2392 -5889 2396 -5884
rect 2399 -5889 2402 -5884
rect 2448 -5889 2452 -5884
rect 2455 -5889 2458 -5884
rect 2509 -5889 2513 -5884
rect 2516 -5889 2519 -5884
rect 2593 -5889 2597 -5884
rect 2600 -5889 2603 -5884
rect 2616 -5889 2620 -5884
rect 2623 -5889 2626 -5884
rect 2639 -5889 2643 -5884
rect 2646 -5889 2649 -5884
rect 2662 -5889 2666 -5884
rect 2669 -5889 2672 -5884
rect 2718 -5889 2722 -5884
rect 2725 -5889 2728 -5884
rect 2783 -5890 2787 -5885
rect 2790 -5890 2793 -5885
rect 2873 -5889 2877 -5884
rect 2880 -5889 2883 -5884
rect 2896 -5889 2900 -5884
rect 2903 -5889 2906 -5884
rect 2919 -5889 2923 -5884
rect 2926 -5889 2929 -5884
rect 2942 -5889 2946 -5884
rect 2949 -5889 2952 -5884
rect 2965 -5889 2969 -5884
rect 2972 -5889 2975 -5884
rect 3021 -5889 3025 -5884
rect 3028 -5889 3031 -5884
rect 2088 -6049 2091 -6045
rect 2094 -6049 2097 -6045
rect 2111 -6049 2114 -6045
rect 2117 -6049 2120 -6045
rect 2141 -6049 2145 -6045
rect 2148 -6049 2151 -6045
rect 2164 -6049 2168 -6045
rect 2171 -6049 2174 -6045
rect 2221 -6027 2225 -6022
rect 2228 -6027 2231 -6022
rect -1577 -6227 -1574 -6223
rect -1571 -6227 -1568 -6223
rect -1554 -6227 -1551 -6223
rect -1548 -6227 -1545 -6223
rect -1524 -6227 -1520 -6223
rect -1517 -6227 -1514 -6223
rect -1501 -6227 -1497 -6223
rect -1494 -6227 -1491 -6223
rect -787 -6227 -784 -6223
rect -781 -6227 -778 -6223
rect -764 -6227 -761 -6223
rect -758 -6227 -755 -6223
rect -734 -6227 -730 -6223
rect -727 -6227 -724 -6223
rect -711 -6227 -707 -6223
rect -704 -6227 -701 -6223
rect 195 -6227 198 -6223
rect 201 -6227 204 -6223
rect 218 -6227 221 -6223
rect 224 -6227 227 -6223
rect 248 -6227 252 -6223
rect 255 -6227 258 -6223
rect 271 -6227 275 -6223
rect 278 -6227 281 -6223
rect 1079 -6227 1082 -6223
rect 1085 -6227 1088 -6223
rect 1102 -6227 1105 -6223
rect 1108 -6227 1111 -6223
rect 1132 -6227 1136 -6223
rect 1139 -6227 1142 -6223
rect 1155 -6227 1159 -6223
rect 1162 -6227 1165 -6223
rect 2087 -6194 2090 -6190
rect 2093 -6194 2096 -6190
rect 2110 -6194 2113 -6190
rect 2116 -6194 2119 -6190
rect 2140 -6194 2144 -6190
rect 2147 -6194 2150 -6190
rect 2163 -6194 2167 -6190
rect 2170 -6194 2173 -6190
rect 2220 -6172 2224 -6167
rect 2227 -6172 2230 -6167
rect 2350 -6264 2354 -6259
rect 2357 -6264 2360 -6259
rect 2373 -6264 2377 -6259
rect 2380 -6264 2383 -6259
rect 2396 -6264 2400 -6259
rect 2403 -6264 2406 -6259
rect 2419 -6264 2423 -6259
rect 2426 -6264 2429 -6259
rect 2475 -6264 2479 -6259
rect 2482 -6264 2485 -6259
rect 2087 -6356 2090 -6352
rect 2093 -6356 2096 -6352
rect 2110 -6356 2113 -6352
rect 2116 -6356 2119 -6352
rect 2140 -6356 2144 -6352
rect 2147 -6356 2150 -6352
rect 2163 -6356 2167 -6352
rect 2170 -6356 2173 -6352
rect 2220 -6334 2224 -6329
rect 2227 -6334 2230 -6329
rect -1564 -6538 -1561 -6534
rect -1558 -6538 -1555 -6534
rect -1541 -6538 -1538 -6534
rect -1535 -6538 -1532 -6534
rect -1511 -6538 -1507 -6534
rect -1504 -6538 -1501 -6534
rect -1488 -6538 -1484 -6534
rect -1481 -6538 -1478 -6534
rect -1409 -6537 -1406 -6533
rect -1403 -6537 -1400 -6533
rect -1386 -6537 -1383 -6533
rect -1380 -6537 -1377 -6533
rect -1356 -6537 -1352 -6533
rect -1349 -6537 -1346 -6533
rect -1333 -6537 -1329 -6533
rect -1326 -6537 -1323 -6533
rect -763 -6536 -760 -6532
rect -757 -6536 -754 -6532
rect -740 -6536 -737 -6532
rect -734 -6536 -731 -6532
rect -710 -6536 -706 -6532
rect -703 -6536 -700 -6532
rect -687 -6536 -683 -6532
rect -680 -6536 -677 -6532
rect -608 -6535 -605 -6531
rect -602 -6535 -599 -6531
rect -585 -6535 -582 -6531
rect -579 -6535 -576 -6531
rect -555 -6535 -551 -6531
rect -548 -6535 -545 -6531
rect -532 -6535 -528 -6531
rect -525 -6535 -522 -6531
rect 140 -6536 143 -6532
rect 146 -6536 149 -6532
rect 163 -6536 166 -6532
rect 169 -6536 172 -6532
rect 193 -6536 197 -6532
rect 200 -6536 203 -6532
rect 216 -6536 220 -6532
rect 223 -6536 226 -6532
rect 295 -6535 298 -6531
rect 301 -6535 304 -6531
rect 318 -6535 321 -6531
rect 324 -6535 327 -6531
rect 348 -6535 352 -6531
rect 355 -6535 358 -6531
rect 371 -6535 375 -6531
rect 378 -6535 381 -6531
rect 1008 -6535 1011 -6531
rect 1014 -6535 1017 -6531
rect 1031 -6535 1034 -6531
rect 1037 -6535 1040 -6531
rect 1061 -6535 1065 -6531
rect 1068 -6535 1071 -6531
rect 1084 -6535 1088 -6531
rect 1091 -6535 1094 -6531
rect 1163 -6534 1166 -6530
rect 1169 -6534 1172 -6530
rect 1186 -6534 1189 -6530
rect 1192 -6534 1195 -6530
rect 1216 -6534 1220 -6530
rect 1223 -6534 1226 -6530
rect 1239 -6534 1243 -6530
rect 1246 -6534 1249 -6530
rect 2088 -6510 2091 -6506
rect 2094 -6510 2097 -6506
rect 2111 -6510 2114 -6506
rect 2117 -6510 2120 -6506
rect 2141 -6510 2145 -6506
rect 2148 -6510 2151 -6506
rect 2164 -6510 2168 -6506
rect 2171 -6510 2174 -6506
rect 2221 -6488 2225 -6483
rect 2228 -6488 2231 -6483
rect -1225 -6665 -1221 -6660
rect -1218 -6665 -1215 -6660
rect -1202 -6665 -1198 -6660
rect -1195 -6665 -1192 -6660
rect -1179 -6665 -1175 -6660
rect -1172 -6665 -1169 -6660
rect -1156 -6665 -1152 -6660
rect -1149 -6665 -1146 -6660
rect -424 -6663 -420 -6658
rect -417 -6663 -414 -6658
rect -401 -6663 -397 -6658
rect -394 -6663 -391 -6658
rect -378 -6663 -374 -6658
rect -371 -6663 -368 -6658
rect -355 -6663 -351 -6658
rect -348 -6663 -345 -6658
rect -1671 -6672 -1667 -6667
rect -1664 -6672 -1661 -6667
rect -1648 -6672 -1644 -6667
rect -1641 -6672 -1638 -6667
rect -1610 -6672 -1606 -6667
rect -1603 -6672 -1600 -6667
rect -1531 -6671 -1527 -6666
rect -1524 -6671 -1521 -6666
rect -1508 -6671 -1504 -6666
rect -1501 -6671 -1498 -6666
rect -1470 -6671 -1466 -6666
rect -1463 -6671 -1460 -6666
rect -1386 -6670 -1382 -6665
rect -1379 -6670 -1376 -6665
rect -1363 -6670 -1359 -6665
rect -1356 -6670 -1353 -6665
rect -1325 -6670 -1321 -6665
rect -1318 -6670 -1315 -6665
rect -870 -6670 -866 -6665
rect -863 -6670 -860 -6665
rect -847 -6670 -843 -6665
rect -840 -6670 -837 -6665
rect -809 -6670 -805 -6665
rect -802 -6670 -799 -6665
rect -730 -6669 -726 -6664
rect -723 -6669 -720 -6664
rect -707 -6669 -703 -6664
rect -700 -6669 -697 -6664
rect -669 -6669 -665 -6664
rect -662 -6669 -659 -6664
rect -585 -6668 -581 -6663
rect -578 -6668 -575 -6663
rect -562 -6668 -558 -6663
rect -555 -6668 -552 -6663
rect -524 -6668 -520 -6663
rect -517 -6668 -514 -6663
rect 479 -6663 483 -6658
rect 486 -6663 489 -6658
rect 502 -6663 506 -6658
rect 509 -6663 512 -6658
rect 525 -6663 529 -6658
rect 532 -6663 535 -6658
rect 548 -6663 552 -6658
rect 555 -6663 558 -6658
rect 33 -6670 37 -6665
rect 40 -6670 43 -6665
rect 56 -6670 60 -6665
rect 63 -6670 66 -6665
rect 94 -6670 98 -6665
rect 101 -6670 104 -6665
rect 173 -6669 177 -6664
rect 180 -6669 183 -6664
rect 196 -6669 200 -6664
rect 203 -6669 206 -6664
rect 234 -6669 238 -6664
rect 241 -6669 244 -6664
rect 318 -6668 322 -6663
rect 325 -6668 328 -6663
rect 341 -6668 345 -6663
rect 348 -6668 351 -6663
rect 379 -6668 383 -6663
rect 386 -6668 389 -6663
rect 1347 -6662 1351 -6657
rect 1354 -6662 1357 -6657
rect 1370 -6662 1374 -6657
rect 1377 -6662 1380 -6657
rect 1393 -6662 1397 -6657
rect 1400 -6662 1403 -6657
rect 1416 -6662 1420 -6657
rect 1423 -6662 1426 -6657
rect 901 -6669 905 -6664
rect 908 -6669 911 -6664
rect 924 -6669 928 -6664
rect 931 -6669 934 -6664
rect 962 -6669 966 -6664
rect 969 -6669 972 -6664
rect 1041 -6668 1045 -6663
rect 1048 -6668 1051 -6663
rect 1064 -6668 1068 -6663
rect 1071 -6668 1074 -6663
rect 1102 -6668 1106 -6663
rect 1109 -6668 1112 -6663
rect 1186 -6667 1190 -6662
rect 1193 -6667 1196 -6662
rect 1209 -6667 1213 -6662
rect 1216 -6667 1219 -6662
rect 1247 -6667 1251 -6662
rect 1254 -6667 1257 -6662
rect 3103 -6682 3107 -6677
rect 3110 -6682 3113 -6677
rect 3126 -6682 3130 -6677
rect 3133 -6682 3136 -6677
rect 3149 -6682 3153 -6677
rect 3156 -6682 3159 -6677
rect 3172 -6682 3176 -6677
rect 3179 -6682 3182 -6677
rect 3195 -6682 3199 -6677
rect 3202 -6682 3205 -6677
rect 2092 -6698 2096 -6693
rect 2099 -6698 2102 -6693
rect 2139 -6697 2143 -6692
rect 2146 -6697 2149 -6692
rect 2162 -6697 2166 -6692
rect 2169 -6697 2172 -6692
rect 2218 -6697 2222 -6692
rect 2225 -6697 2228 -6692
rect 2283 -6697 2287 -6692
rect 2290 -6697 2293 -6692
rect 2348 -6697 2352 -6692
rect 2355 -6697 2358 -6692
rect 2371 -6697 2375 -6692
rect 2378 -6697 2381 -6692
rect 2394 -6697 2398 -6692
rect 2401 -6697 2404 -6692
rect 2450 -6697 2454 -6692
rect 2457 -6697 2460 -6692
rect 2510 -6697 2514 -6692
rect 2517 -6697 2520 -6692
rect 2594 -6697 2598 -6692
rect 2601 -6697 2604 -6692
rect 2617 -6697 2621 -6692
rect 2624 -6697 2627 -6692
rect 2640 -6697 2644 -6692
rect 2647 -6697 2650 -6692
rect 2663 -6697 2667 -6692
rect 2670 -6697 2673 -6692
rect 2719 -6697 2723 -6692
rect 2726 -6697 2729 -6692
rect 2781 -6697 2785 -6692
rect 2788 -6697 2791 -6692
rect 2871 -6696 2875 -6691
rect 2878 -6696 2881 -6691
rect 2894 -6696 2898 -6691
rect 2901 -6696 2904 -6691
rect 2917 -6696 2921 -6691
rect 2924 -6696 2927 -6691
rect 2940 -6696 2944 -6691
rect 2947 -6696 2950 -6691
rect 2963 -6696 2967 -6691
rect 2970 -6696 2973 -6691
rect 3019 -6696 3023 -6691
rect 3026 -6696 3029 -6691
<< pdiffusion >>
rect 666 -5016 669 -5010
rect 672 -5016 675 -5010
rect 689 -5016 692 -5010
rect 695 -5016 698 -5010
rect 727 -5016 730 -5010
rect 733 -5016 736 -5010
rect 1118 -5101 1121 -5095
rect 1124 -5101 1127 -5095
rect 970 -5118 973 -5112
rect 976 -5118 979 -5112
rect 993 -5118 996 -5112
rect 999 -5118 1002 -5112
rect 1031 -5118 1034 -5112
rect 1037 -5118 1040 -5112
rect 1208 -5114 1211 -5108
rect 1214 -5114 1217 -5108
rect 1231 -5114 1234 -5108
rect 1237 -5114 1240 -5108
rect 1269 -5114 1272 -5108
rect 1275 -5114 1278 -5108
rect 1339 -5114 1342 -5108
rect 1345 -5114 1348 -5108
rect 1362 -5114 1365 -5108
rect 1368 -5114 1371 -5108
rect 1400 -5114 1403 -5108
rect 1406 -5114 1409 -5108
rect 1495 -5114 1498 -5108
rect 1501 -5114 1504 -5108
rect 1518 -5114 1521 -5108
rect 1524 -5114 1527 -5108
rect 1556 -5114 1559 -5108
rect 1562 -5114 1565 -5108
rect 1117 -5169 1120 -5163
rect 1123 -5169 1126 -5163
rect 572 -5326 575 -5320
rect 578 -5326 581 -5320
rect 595 -5326 598 -5320
rect 601 -5326 604 -5320
rect 638 -5326 641 -5320
rect 644 -5326 647 -5320
rect 680 -5326 683 -5320
rect 686 -5326 689 -5320
rect 703 -5326 706 -5320
rect 709 -5326 712 -5320
rect 746 -5326 749 -5320
rect 752 -5326 755 -5320
rect 792 -5326 795 -5320
rect 798 -5326 801 -5320
rect 815 -5326 818 -5320
rect 821 -5326 824 -5320
rect 858 -5326 861 -5320
rect 864 -5326 867 -5320
rect 904 -5326 907 -5320
rect 910 -5326 913 -5320
rect 927 -5326 930 -5320
rect 933 -5326 936 -5320
rect 970 -5326 973 -5320
rect 976 -5326 979 -5320
rect 1015 -5326 1018 -5320
rect 1021 -5326 1024 -5320
rect 1038 -5326 1041 -5320
rect 1044 -5326 1047 -5320
rect 1081 -5326 1084 -5320
rect 1087 -5326 1090 -5320
rect 1127 -5326 1130 -5320
rect 1133 -5326 1136 -5320
rect 1150 -5326 1153 -5320
rect 1156 -5326 1159 -5320
rect 1193 -5326 1196 -5320
rect 1199 -5326 1202 -5320
rect 1239 -5326 1242 -5320
rect 1245 -5326 1248 -5320
rect 1262 -5326 1265 -5320
rect 1268 -5326 1271 -5320
rect 1305 -5326 1308 -5320
rect 1311 -5326 1314 -5320
rect 1351 -5326 1354 -5320
rect 1357 -5326 1360 -5320
rect 1374 -5326 1377 -5320
rect 1380 -5326 1383 -5320
rect 1417 -5326 1420 -5320
rect 1423 -5326 1426 -5320
rect 1791 -5324 1794 -5318
rect 1797 -5324 1800 -5318
rect 1814 -5324 1817 -5318
rect 1820 -5324 1823 -5318
rect 1857 -5324 1860 -5318
rect 1863 -5324 1866 -5318
rect 1899 -5324 1902 -5318
rect 1905 -5324 1908 -5318
rect 1922 -5324 1925 -5318
rect 1928 -5324 1931 -5318
rect 1965 -5324 1968 -5318
rect 1971 -5324 1974 -5318
rect 2011 -5324 2014 -5318
rect 2017 -5324 2020 -5318
rect 2034 -5324 2037 -5318
rect 2040 -5324 2043 -5318
rect 2077 -5324 2080 -5318
rect 2083 -5324 2086 -5318
rect 2123 -5324 2126 -5318
rect 2129 -5324 2132 -5318
rect 2146 -5324 2149 -5318
rect 2152 -5324 2155 -5318
rect 2189 -5324 2192 -5318
rect 2195 -5324 2198 -5318
rect 2234 -5324 2237 -5318
rect 2240 -5324 2243 -5318
rect 2257 -5324 2260 -5318
rect 2263 -5324 2266 -5318
rect 2300 -5324 2303 -5318
rect 2306 -5324 2309 -5318
rect 2346 -5324 2349 -5318
rect 2352 -5324 2355 -5318
rect 2369 -5324 2372 -5318
rect 2375 -5324 2378 -5318
rect 2412 -5324 2415 -5318
rect 2418 -5324 2421 -5318
rect 2458 -5324 2461 -5318
rect 2464 -5324 2467 -5318
rect 2481 -5324 2484 -5318
rect 2487 -5324 2490 -5318
rect 2524 -5324 2527 -5318
rect 2530 -5324 2533 -5318
rect 2570 -5324 2573 -5318
rect 2576 -5324 2579 -5318
rect 2593 -5324 2596 -5318
rect 2599 -5324 2602 -5318
rect 2636 -5324 2639 -5318
rect 2642 -5324 2645 -5318
rect -579 -5333 -576 -5327
rect -573 -5333 -570 -5327
rect -556 -5333 -553 -5327
rect -550 -5333 -547 -5327
rect -513 -5333 -510 -5327
rect -507 -5333 -504 -5327
rect -471 -5333 -468 -5327
rect -465 -5333 -462 -5327
rect -448 -5333 -445 -5327
rect -442 -5333 -439 -5327
rect -405 -5333 -402 -5327
rect -399 -5333 -396 -5327
rect -359 -5333 -356 -5327
rect -353 -5333 -350 -5327
rect -336 -5333 -333 -5327
rect -330 -5333 -327 -5327
rect -293 -5333 -290 -5327
rect -287 -5333 -284 -5327
rect -247 -5333 -244 -5327
rect -241 -5333 -238 -5327
rect -224 -5333 -221 -5327
rect -218 -5333 -215 -5327
rect -181 -5333 -178 -5327
rect -175 -5333 -172 -5327
rect -136 -5333 -133 -5327
rect -130 -5333 -127 -5327
rect -113 -5333 -110 -5327
rect -107 -5333 -104 -5327
rect -70 -5333 -67 -5327
rect -64 -5333 -61 -5327
rect -24 -5333 -21 -5327
rect -18 -5333 -15 -5327
rect -1 -5333 2 -5327
rect 5 -5333 8 -5327
rect 42 -5333 45 -5327
rect 48 -5333 51 -5327
rect 88 -5333 91 -5327
rect 94 -5333 97 -5327
rect 111 -5333 114 -5327
rect 117 -5333 120 -5327
rect 154 -5333 157 -5327
rect 160 -5333 163 -5327
rect 200 -5333 203 -5327
rect 206 -5333 209 -5327
rect 223 -5333 226 -5327
rect 229 -5333 232 -5327
rect 266 -5333 269 -5327
rect 272 -5333 275 -5327
rect 2574 -5715 2577 -5709
rect 2580 -5715 2583 -5709
rect 2597 -5715 2600 -5709
rect 2603 -5715 2606 -5709
rect 2620 -5715 2623 -5709
rect 2626 -5715 2629 -5709
rect 2643 -5715 2646 -5709
rect 2649 -5715 2652 -5709
rect 2666 -5715 2669 -5709
rect 2672 -5715 2675 -5709
rect -545 -5817 -542 -5811
rect -539 -5817 -536 -5811
rect -522 -5817 -519 -5811
rect -516 -5817 -513 -5811
rect -484 -5817 -481 -5811
rect -478 -5817 -475 -5811
rect -406 -5817 -403 -5811
rect -400 -5817 -397 -5811
rect -383 -5817 -380 -5811
rect -377 -5817 -374 -5811
rect -345 -5817 -342 -5811
rect -339 -5817 -336 -5811
rect -268 -5817 -265 -5811
rect -262 -5817 -259 -5811
rect -245 -5817 -242 -5811
rect -239 -5817 -236 -5811
rect -207 -5817 -204 -5811
rect -201 -5817 -198 -5811
rect -118 -5817 -115 -5811
rect -112 -5817 -109 -5811
rect -95 -5817 -92 -5811
rect -89 -5817 -86 -5811
rect -57 -5817 -54 -5811
rect -51 -5817 -48 -5811
rect 2146 -5853 2149 -5847
rect 2152 -5853 2155 -5847
rect 2169 -5853 2172 -5847
rect 2175 -5853 2178 -5847
rect 2225 -5853 2228 -5847
rect 2231 -5853 2234 -5847
rect 2347 -5853 2350 -5847
rect 2353 -5853 2356 -5847
rect 2370 -5853 2373 -5847
rect 2376 -5853 2379 -5847
rect 2393 -5853 2396 -5847
rect 2399 -5853 2402 -5847
rect 2449 -5853 2452 -5847
rect 2455 -5853 2458 -5847
rect 2594 -5853 2597 -5847
rect 2600 -5853 2603 -5847
rect 2617 -5853 2620 -5847
rect 2623 -5853 2626 -5847
rect 2640 -5853 2643 -5847
rect 2646 -5853 2649 -5847
rect 2663 -5853 2666 -5847
rect 2669 -5853 2672 -5847
rect 2719 -5853 2722 -5847
rect 2725 -5853 2728 -5847
rect 2874 -5853 2877 -5847
rect 2880 -5853 2883 -5847
rect 2897 -5853 2900 -5847
rect 2903 -5853 2906 -5847
rect 2920 -5853 2923 -5847
rect 2926 -5853 2929 -5847
rect 2943 -5853 2946 -5847
rect 2949 -5853 2952 -5847
rect 2966 -5853 2969 -5847
rect 2972 -5853 2975 -5847
rect 3022 -5853 3025 -5847
rect 3028 -5853 3031 -5847
rect 2099 -5864 2102 -5858
rect 2105 -5864 2108 -5858
rect 2282 -5863 2285 -5857
rect 2288 -5863 2291 -5857
rect 2510 -5863 2513 -5857
rect 2516 -5863 2519 -5857
rect 2784 -5864 2787 -5858
rect 2790 -5864 2793 -5858
rect 2088 -5996 2091 -5990
rect 2094 -5996 2097 -5990
rect 2111 -5996 2114 -5990
rect 2117 -5996 2120 -5990
rect 2142 -5996 2145 -5990
rect 2148 -5996 2151 -5990
rect 2165 -5996 2168 -5990
rect 2171 -5996 2174 -5990
rect 2222 -6001 2225 -5995
rect 2228 -6001 2231 -5995
rect -1577 -6174 -1574 -6168
rect -1571 -6174 -1568 -6168
rect -1554 -6174 -1551 -6168
rect -1548 -6174 -1545 -6168
rect -1523 -6174 -1520 -6168
rect -1517 -6174 -1514 -6168
rect -1500 -6174 -1497 -6168
rect -1494 -6174 -1491 -6168
rect -787 -6174 -784 -6168
rect -781 -6174 -778 -6168
rect -764 -6174 -761 -6168
rect -758 -6174 -755 -6168
rect -733 -6174 -730 -6168
rect -727 -6174 -724 -6168
rect -710 -6174 -707 -6168
rect -704 -6174 -701 -6168
rect 195 -6174 198 -6168
rect 201 -6174 204 -6168
rect 218 -6174 221 -6168
rect 224 -6174 227 -6168
rect 249 -6174 252 -6168
rect 255 -6174 258 -6168
rect 272 -6174 275 -6168
rect 278 -6174 281 -6168
rect 1079 -6174 1082 -6168
rect 1085 -6174 1088 -6168
rect 1102 -6174 1105 -6168
rect 1108 -6174 1111 -6168
rect 1133 -6174 1136 -6168
rect 1139 -6174 1142 -6168
rect 1156 -6174 1159 -6168
rect 1162 -6174 1165 -6168
rect 2087 -6141 2090 -6135
rect 2093 -6141 2096 -6135
rect 2110 -6141 2113 -6135
rect 2116 -6141 2119 -6135
rect 2141 -6141 2144 -6135
rect 2147 -6141 2150 -6135
rect 2164 -6141 2167 -6135
rect 2170 -6141 2173 -6135
rect 2221 -6146 2224 -6140
rect 2227 -6146 2230 -6140
rect 2351 -6228 2354 -6222
rect 2357 -6228 2360 -6222
rect 2374 -6228 2377 -6222
rect 2380 -6228 2383 -6222
rect 2397 -6228 2400 -6222
rect 2403 -6228 2406 -6222
rect 2420 -6228 2423 -6222
rect 2426 -6228 2429 -6222
rect 2476 -6228 2479 -6222
rect 2482 -6228 2485 -6222
rect 2087 -6303 2090 -6297
rect 2093 -6303 2096 -6297
rect 2110 -6303 2113 -6297
rect 2116 -6303 2119 -6297
rect 2141 -6303 2144 -6297
rect 2147 -6303 2150 -6297
rect 2164 -6303 2167 -6297
rect 2170 -6303 2173 -6297
rect 2221 -6308 2224 -6302
rect 2227 -6308 2230 -6302
rect -1564 -6485 -1561 -6479
rect -1558 -6485 -1555 -6479
rect -1541 -6485 -1538 -6479
rect -1535 -6485 -1532 -6479
rect -1510 -6485 -1507 -6479
rect -1504 -6485 -1501 -6479
rect -1487 -6485 -1484 -6479
rect -1481 -6485 -1478 -6479
rect -1409 -6484 -1406 -6478
rect -1403 -6484 -1400 -6478
rect -1386 -6484 -1383 -6478
rect -1380 -6484 -1377 -6478
rect -1355 -6484 -1352 -6478
rect -1349 -6484 -1346 -6478
rect -1332 -6484 -1329 -6478
rect -1326 -6484 -1323 -6478
rect -763 -6483 -760 -6477
rect -757 -6483 -754 -6477
rect -740 -6483 -737 -6477
rect -734 -6483 -731 -6477
rect -709 -6483 -706 -6477
rect -703 -6483 -700 -6477
rect -686 -6483 -683 -6477
rect -680 -6483 -677 -6477
rect -608 -6482 -605 -6476
rect -602 -6482 -599 -6476
rect -585 -6482 -582 -6476
rect -579 -6482 -576 -6476
rect -554 -6482 -551 -6476
rect -548 -6482 -545 -6476
rect -531 -6482 -528 -6476
rect -525 -6482 -522 -6476
rect 140 -6483 143 -6477
rect 146 -6483 149 -6477
rect 163 -6483 166 -6477
rect 169 -6483 172 -6477
rect 194 -6483 197 -6477
rect 200 -6483 203 -6477
rect 217 -6483 220 -6477
rect 223 -6483 226 -6477
rect 295 -6482 298 -6476
rect 301 -6482 304 -6476
rect 318 -6482 321 -6476
rect 324 -6482 327 -6476
rect 349 -6482 352 -6476
rect 355 -6482 358 -6476
rect 372 -6482 375 -6476
rect 378 -6482 381 -6476
rect 1008 -6482 1011 -6476
rect 1014 -6482 1017 -6476
rect 1031 -6482 1034 -6476
rect 1037 -6482 1040 -6476
rect 1062 -6482 1065 -6476
rect 1068 -6482 1071 -6476
rect 1085 -6482 1088 -6476
rect 1091 -6482 1094 -6476
rect 1163 -6481 1166 -6475
rect 1169 -6481 1172 -6475
rect 1186 -6481 1189 -6475
rect 1192 -6481 1195 -6475
rect 1217 -6481 1220 -6475
rect 1223 -6481 1226 -6475
rect 1240 -6481 1243 -6475
rect 1246 -6481 1249 -6475
rect 2088 -6457 2091 -6451
rect 2094 -6457 2097 -6451
rect 2111 -6457 2114 -6451
rect 2117 -6457 2120 -6451
rect 2142 -6457 2145 -6451
rect 2148 -6457 2151 -6451
rect 2165 -6457 2168 -6451
rect 2171 -6457 2174 -6451
rect 2222 -6462 2225 -6456
rect 2228 -6462 2231 -6456
rect -1670 -6636 -1667 -6630
rect -1664 -6636 -1661 -6630
rect -1647 -6636 -1644 -6630
rect -1641 -6636 -1638 -6630
rect -1609 -6636 -1606 -6630
rect -1603 -6636 -1600 -6630
rect -1530 -6635 -1527 -6629
rect -1524 -6635 -1521 -6629
rect -1507 -6635 -1504 -6629
rect -1501 -6635 -1498 -6629
rect -1469 -6635 -1466 -6629
rect -1463 -6635 -1460 -6629
rect -1385 -6634 -1382 -6628
rect -1379 -6634 -1376 -6628
rect -1362 -6634 -1359 -6628
rect -1356 -6634 -1353 -6628
rect -1324 -6634 -1321 -6628
rect -1318 -6634 -1315 -6628
rect -1224 -6637 -1221 -6631
rect -1218 -6637 -1215 -6631
rect -1201 -6637 -1198 -6631
rect -1195 -6637 -1192 -6631
rect -1178 -6637 -1175 -6631
rect -1172 -6637 -1169 -6631
rect -1155 -6637 -1152 -6631
rect -1149 -6637 -1146 -6631
rect -869 -6634 -866 -6628
rect -863 -6634 -860 -6628
rect -846 -6634 -843 -6628
rect -840 -6634 -837 -6628
rect -808 -6634 -805 -6628
rect -802 -6634 -799 -6628
rect -729 -6633 -726 -6627
rect -723 -6633 -720 -6627
rect -706 -6633 -703 -6627
rect -700 -6633 -697 -6627
rect -668 -6633 -665 -6627
rect -662 -6633 -659 -6627
rect -584 -6632 -581 -6626
rect -578 -6632 -575 -6626
rect -561 -6632 -558 -6626
rect -555 -6632 -552 -6626
rect -523 -6632 -520 -6626
rect -517 -6632 -514 -6626
rect -423 -6635 -420 -6629
rect -417 -6635 -414 -6629
rect -400 -6635 -397 -6629
rect -394 -6635 -391 -6629
rect -377 -6635 -374 -6629
rect -371 -6635 -368 -6629
rect -354 -6635 -351 -6629
rect -348 -6635 -345 -6629
rect 34 -6634 37 -6628
rect 40 -6634 43 -6628
rect 57 -6634 60 -6628
rect 63 -6634 66 -6628
rect 95 -6634 98 -6628
rect 101 -6634 104 -6628
rect 174 -6633 177 -6627
rect 180 -6633 183 -6627
rect 197 -6633 200 -6627
rect 203 -6633 206 -6627
rect 235 -6633 238 -6627
rect 241 -6633 244 -6627
rect 319 -6632 322 -6626
rect 325 -6632 328 -6626
rect 342 -6632 345 -6626
rect 348 -6632 351 -6626
rect 380 -6632 383 -6626
rect 386 -6632 389 -6626
rect 480 -6635 483 -6629
rect 486 -6635 489 -6629
rect 503 -6635 506 -6629
rect 509 -6635 512 -6629
rect 526 -6635 529 -6629
rect 532 -6635 535 -6629
rect 549 -6635 552 -6629
rect 555 -6635 558 -6629
rect 902 -6633 905 -6627
rect 908 -6633 911 -6627
rect 925 -6633 928 -6627
rect 931 -6633 934 -6627
rect 963 -6633 966 -6627
rect 969 -6633 972 -6627
rect 1042 -6632 1045 -6626
rect 1048 -6632 1051 -6626
rect 1065 -6632 1068 -6626
rect 1071 -6632 1074 -6626
rect 1103 -6632 1106 -6626
rect 1109 -6632 1112 -6626
rect 1187 -6631 1190 -6625
rect 1193 -6631 1196 -6625
rect 1210 -6631 1213 -6625
rect 1216 -6631 1219 -6625
rect 1248 -6631 1251 -6625
rect 1254 -6631 1257 -6625
rect 1348 -6634 1351 -6628
rect 1354 -6634 1357 -6628
rect 1371 -6634 1374 -6628
rect 1377 -6634 1380 -6628
rect 1394 -6634 1397 -6628
rect 1400 -6634 1403 -6628
rect 1417 -6634 1420 -6628
rect 1423 -6634 1426 -6628
rect 3104 -6654 3107 -6648
rect 3110 -6654 3113 -6648
rect 3127 -6654 3130 -6648
rect 3133 -6654 3136 -6648
rect 3150 -6654 3153 -6648
rect 3156 -6654 3159 -6648
rect 3173 -6654 3176 -6648
rect 3179 -6654 3182 -6648
rect 3196 -6654 3199 -6648
rect 3202 -6654 3205 -6648
rect 2140 -6661 2143 -6655
rect 2146 -6661 2149 -6655
rect 2163 -6661 2166 -6655
rect 2169 -6661 2172 -6655
rect 2219 -6661 2222 -6655
rect 2225 -6661 2228 -6655
rect 2349 -6661 2352 -6655
rect 2355 -6661 2358 -6655
rect 2372 -6661 2375 -6655
rect 2378 -6661 2381 -6655
rect 2395 -6661 2398 -6655
rect 2401 -6661 2404 -6655
rect 2451 -6661 2454 -6655
rect 2457 -6661 2460 -6655
rect 2595 -6661 2598 -6655
rect 2601 -6661 2604 -6655
rect 2618 -6661 2621 -6655
rect 2624 -6661 2627 -6655
rect 2641 -6661 2644 -6655
rect 2647 -6661 2650 -6655
rect 2664 -6661 2667 -6655
rect 2670 -6661 2673 -6655
rect 2720 -6661 2723 -6655
rect 2726 -6661 2729 -6655
rect 2872 -6660 2875 -6654
rect 2878 -6660 2881 -6654
rect 2895 -6660 2898 -6654
rect 2901 -6660 2904 -6654
rect 2918 -6660 2921 -6654
rect 2924 -6660 2927 -6654
rect 2941 -6660 2944 -6654
rect 2947 -6660 2950 -6654
rect 2964 -6660 2967 -6654
rect 2970 -6660 2973 -6654
rect 3020 -6660 3023 -6654
rect 3026 -6660 3029 -6654
rect 2093 -6672 2096 -6666
rect 2099 -6672 2102 -6666
rect 2284 -6671 2287 -6665
rect 2290 -6671 2293 -6665
rect 2511 -6671 2514 -6665
rect 2517 -6671 2520 -6665
rect 2782 -6671 2785 -6665
rect 2788 -6671 2791 -6665
<< ndcontact >>
rect 661 -5052 665 -5047
rect 675 -5052 679 -5047
rect 684 -5052 688 -5047
rect 698 -5052 702 -5047
rect 722 -5052 726 -5047
rect 736 -5052 740 -5047
rect 1113 -5127 1117 -5122
rect 1127 -5127 1131 -5122
rect 965 -5154 969 -5149
rect 979 -5154 983 -5149
rect 988 -5154 992 -5149
rect 1002 -5154 1006 -5149
rect 1026 -5154 1030 -5149
rect 1040 -5154 1044 -5149
rect 1203 -5150 1207 -5145
rect 1217 -5150 1221 -5145
rect 1226 -5150 1230 -5145
rect 1240 -5150 1244 -5145
rect 1264 -5150 1268 -5145
rect 1278 -5150 1282 -5145
rect 1334 -5150 1338 -5145
rect 1348 -5150 1352 -5145
rect 1357 -5150 1361 -5145
rect 1371 -5150 1375 -5145
rect 1395 -5150 1399 -5145
rect 1409 -5150 1413 -5145
rect 1490 -5150 1494 -5145
rect 1504 -5150 1508 -5145
rect 1513 -5150 1517 -5145
rect 1527 -5150 1531 -5145
rect 1551 -5150 1555 -5145
rect 1565 -5150 1569 -5145
rect 1112 -5195 1116 -5190
rect 1126 -5195 1130 -5190
rect 567 -5362 571 -5357
rect 581 -5362 585 -5357
rect 590 -5362 594 -5357
rect 604 -5362 608 -5357
rect 633 -5362 637 -5357
rect 647 -5362 651 -5357
rect 675 -5362 679 -5357
rect 689 -5362 693 -5357
rect 698 -5362 702 -5357
rect 712 -5362 716 -5357
rect 741 -5362 745 -5357
rect 755 -5362 759 -5357
rect 787 -5362 791 -5357
rect 801 -5362 805 -5357
rect 810 -5362 814 -5357
rect 824 -5362 828 -5357
rect 853 -5362 857 -5357
rect 867 -5362 871 -5357
rect 899 -5362 903 -5357
rect 913 -5362 917 -5357
rect 922 -5362 926 -5357
rect 936 -5362 940 -5357
rect 965 -5362 969 -5357
rect 979 -5362 983 -5357
rect 1010 -5362 1014 -5357
rect 1024 -5362 1028 -5357
rect 1033 -5362 1037 -5357
rect 1047 -5362 1051 -5357
rect 1076 -5362 1080 -5357
rect 1090 -5362 1094 -5357
rect 1122 -5362 1126 -5357
rect 1136 -5362 1140 -5357
rect 1145 -5362 1149 -5357
rect 1159 -5362 1163 -5357
rect 1188 -5362 1192 -5357
rect 1202 -5362 1206 -5357
rect 1234 -5362 1238 -5357
rect 1248 -5362 1252 -5357
rect 1257 -5362 1261 -5357
rect 1271 -5362 1275 -5357
rect 1300 -5362 1304 -5357
rect 1314 -5362 1318 -5357
rect 1346 -5362 1350 -5357
rect 1360 -5362 1364 -5357
rect 1369 -5362 1373 -5357
rect 1383 -5362 1387 -5357
rect 1412 -5362 1416 -5357
rect 1426 -5362 1430 -5357
rect 1786 -5360 1790 -5355
rect 1800 -5360 1804 -5355
rect 1809 -5360 1813 -5355
rect 1823 -5360 1827 -5355
rect 1852 -5360 1856 -5355
rect 1866 -5360 1870 -5355
rect 1894 -5360 1898 -5355
rect 1908 -5360 1912 -5355
rect 1917 -5360 1921 -5355
rect 1931 -5360 1935 -5355
rect 1960 -5360 1964 -5355
rect 1974 -5360 1978 -5355
rect 2006 -5360 2010 -5355
rect 2020 -5360 2024 -5355
rect 2029 -5360 2033 -5355
rect 2043 -5360 2047 -5355
rect 2072 -5360 2076 -5355
rect 2086 -5360 2090 -5355
rect 2118 -5360 2122 -5355
rect 2132 -5360 2136 -5355
rect 2141 -5360 2145 -5355
rect 2155 -5360 2159 -5355
rect 2184 -5360 2188 -5355
rect 2198 -5360 2202 -5355
rect 2229 -5360 2233 -5355
rect 2243 -5360 2247 -5355
rect 2252 -5360 2256 -5355
rect 2266 -5360 2270 -5355
rect 2295 -5360 2299 -5355
rect 2309 -5360 2313 -5355
rect 2341 -5360 2345 -5355
rect 2355 -5360 2359 -5355
rect 2364 -5360 2368 -5355
rect 2378 -5360 2382 -5355
rect 2407 -5360 2411 -5355
rect 2421 -5360 2425 -5355
rect 2453 -5360 2457 -5355
rect 2467 -5360 2471 -5355
rect 2476 -5360 2480 -5355
rect 2490 -5360 2494 -5355
rect 2519 -5360 2523 -5355
rect 2533 -5360 2537 -5355
rect 2565 -5360 2569 -5355
rect 2579 -5360 2583 -5355
rect 2588 -5360 2592 -5355
rect 2602 -5360 2606 -5355
rect 2631 -5360 2635 -5355
rect 2645 -5360 2649 -5355
rect -584 -5369 -580 -5364
rect -570 -5369 -566 -5364
rect -561 -5369 -557 -5364
rect -547 -5369 -543 -5364
rect -518 -5369 -514 -5364
rect -504 -5369 -500 -5364
rect -476 -5369 -472 -5364
rect -462 -5369 -458 -5364
rect -453 -5369 -449 -5364
rect -439 -5369 -435 -5364
rect -410 -5369 -406 -5364
rect -396 -5369 -392 -5364
rect -364 -5369 -360 -5364
rect -350 -5369 -346 -5364
rect -341 -5369 -337 -5364
rect -327 -5369 -323 -5364
rect -298 -5369 -294 -5364
rect -284 -5369 -280 -5364
rect -252 -5369 -248 -5364
rect -238 -5369 -234 -5364
rect -229 -5369 -225 -5364
rect -215 -5369 -211 -5364
rect -186 -5369 -182 -5364
rect -172 -5369 -168 -5364
rect -141 -5369 -137 -5364
rect -127 -5369 -123 -5364
rect -118 -5369 -114 -5364
rect -104 -5369 -100 -5364
rect -75 -5369 -71 -5364
rect -61 -5369 -57 -5364
rect -29 -5369 -25 -5364
rect -15 -5369 -11 -5364
rect -6 -5369 -2 -5364
rect 8 -5369 12 -5364
rect 37 -5369 41 -5364
rect 51 -5369 55 -5364
rect 83 -5369 87 -5364
rect 97 -5369 101 -5364
rect 106 -5369 110 -5364
rect 120 -5369 124 -5364
rect 149 -5369 153 -5364
rect 163 -5369 167 -5364
rect 195 -5369 199 -5364
rect 209 -5369 213 -5364
rect 218 -5369 222 -5364
rect 232 -5369 236 -5364
rect 261 -5369 265 -5364
rect 275 -5369 279 -5364
rect 2569 -5743 2573 -5738
rect 2583 -5743 2587 -5738
rect 2592 -5743 2596 -5738
rect 2606 -5743 2610 -5738
rect 2615 -5743 2619 -5738
rect 2629 -5743 2633 -5738
rect 2638 -5743 2642 -5738
rect 2652 -5743 2656 -5738
rect 2661 -5743 2665 -5738
rect 2675 -5743 2679 -5738
rect -550 -5853 -546 -5848
rect -536 -5853 -532 -5848
rect -527 -5853 -523 -5848
rect -513 -5853 -509 -5848
rect -489 -5853 -485 -5848
rect -475 -5853 -471 -5848
rect -411 -5853 -407 -5848
rect -397 -5853 -393 -5848
rect -388 -5853 -384 -5848
rect -374 -5853 -370 -5848
rect -350 -5853 -346 -5848
rect -336 -5853 -332 -5848
rect -273 -5853 -269 -5848
rect -259 -5853 -255 -5848
rect -250 -5853 -246 -5848
rect -236 -5853 -232 -5848
rect -212 -5853 -208 -5848
rect -198 -5853 -194 -5848
rect -123 -5853 -119 -5848
rect -109 -5853 -105 -5848
rect -100 -5853 -96 -5848
rect -86 -5853 -82 -5848
rect -62 -5853 -58 -5848
rect -48 -5853 -44 -5848
rect 2094 -5890 2098 -5885
rect 2108 -5890 2112 -5885
rect 2141 -5889 2145 -5884
rect 2155 -5889 2159 -5884
rect 2164 -5889 2168 -5884
rect 2178 -5889 2182 -5884
rect 2220 -5889 2224 -5884
rect 2234 -5889 2238 -5884
rect 2277 -5889 2281 -5884
rect 2291 -5889 2295 -5884
rect 2342 -5889 2346 -5884
rect 2356 -5889 2360 -5884
rect 2365 -5889 2369 -5884
rect 2379 -5889 2383 -5884
rect 2388 -5889 2392 -5884
rect 2402 -5889 2406 -5884
rect 2444 -5889 2448 -5884
rect 2458 -5889 2462 -5884
rect 2505 -5889 2509 -5884
rect 2519 -5889 2523 -5884
rect 2589 -5889 2593 -5884
rect 2603 -5889 2607 -5884
rect 2612 -5889 2616 -5884
rect 2626 -5889 2630 -5884
rect 2635 -5889 2639 -5884
rect 2649 -5889 2653 -5884
rect 2658 -5889 2662 -5884
rect 2672 -5889 2676 -5884
rect 2714 -5889 2718 -5884
rect 2728 -5889 2732 -5884
rect 2779 -5890 2783 -5885
rect 2793 -5890 2797 -5885
rect 2869 -5889 2873 -5884
rect 2883 -5889 2887 -5884
rect 2892 -5889 2896 -5884
rect 2906 -5889 2910 -5884
rect 2915 -5889 2919 -5884
rect 2929 -5889 2933 -5884
rect 2938 -5889 2942 -5884
rect 2952 -5889 2956 -5884
rect 2961 -5889 2965 -5884
rect 2975 -5889 2979 -5884
rect 3017 -5889 3021 -5884
rect 3031 -5889 3035 -5884
rect 2083 -6049 2088 -6045
rect 2097 -6049 2101 -6045
rect 2106 -6049 2111 -6045
rect 2120 -6049 2124 -6045
rect 2137 -6049 2141 -6045
rect 2151 -6049 2155 -6045
rect 2160 -6049 2164 -6045
rect 2174 -6049 2178 -6045
rect 2217 -6027 2221 -6022
rect 2231 -6027 2235 -6022
rect -1582 -6227 -1577 -6223
rect -1568 -6227 -1564 -6223
rect -1559 -6227 -1554 -6223
rect -1545 -6227 -1541 -6223
rect -1528 -6227 -1524 -6223
rect -1514 -6227 -1510 -6223
rect -1505 -6227 -1501 -6223
rect -1491 -6227 -1487 -6223
rect -792 -6227 -787 -6223
rect -778 -6227 -774 -6223
rect -769 -6227 -764 -6223
rect -755 -6227 -751 -6223
rect -738 -6227 -734 -6223
rect -724 -6227 -720 -6223
rect -715 -6227 -711 -6223
rect -701 -6227 -697 -6223
rect 190 -6227 195 -6223
rect 204 -6227 208 -6223
rect 213 -6227 218 -6223
rect 227 -6227 231 -6223
rect 244 -6227 248 -6223
rect 258 -6227 262 -6223
rect 267 -6227 271 -6223
rect 281 -6227 285 -6223
rect 1074 -6227 1079 -6223
rect 1088 -6227 1092 -6223
rect 1097 -6227 1102 -6223
rect 1111 -6227 1115 -6223
rect 1128 -6227 1132 -6223
rect 1142 -6227 1146 -6223
rect 1151 -6227 1155 -6223
rect 1165 -6227 1169 -6223
rect 2082 -6194 2087 -6190
rect 2096 -6194 2100 -6190
rect 2105 -6194 2110 -6190
rect 2119 -6194 2123 -6190
rect 2136 -6194 2140 -6190
rect 2150 -6194 2154 -6190
rect 2159 -6194 2163 -6190
rect 2173 -6194 2177 -6190
rect 2216 -6172 2220 -6167
rect 2230 -6172 2234 -6167
rect 2346 -6264 2350 -6259
rect 2360 -6264 2364 -6259
rect 2369 -6264 2373 -6259
rect 2383 -6264 2387 -6259
rect 2392 -6264 2396 -6259
rect 2406 -6264 2410 -6259
rect 2415 -6264 2419 -6259
rect 2429 -6264 2433 -6259
rect 2471 -6264 2475 -6259
rect 2485 -6264 2489 -6259
rect 2082 -6356 2087 -6352
rect 2096 -6356 2100 -6352
rect 2105 -6356 2110 -6352
rect 2119 -6356 2123 -6352
rect 2136 -6356 2140 -6352
rect 2150 -6356 2154 -6352
rect 2159 -6356 2163 -6352
rect 2173 -6356 2177 -6352
rect 2216 -6334 2220 -6329
rect 2230 -6334 2234 -6329
rect -1569 -6538 -1564 -6534
rect -1555 -6538 -1551 -6534
rect -1546 -6538 -1541 -6534
rect -1532 -6538 -1528 -6534
rect -1515 -6538 -1511 -6534
rect -1501 -6538 -1497 -6534
rect -1492 -6538 -1488 -6534
rect -1478 -6538 -1474 -6534
rect -1414 -6537 -1409 -6533
rect -1400 -6537 -1396 -6533
rect -1391 -6537 -1386 -6533
rect -1377 -6537 -1373 -6533
rect -1360 -6537 -1356 -6533
rect -1346 -6537 -1342 -6533
rect -1337 -6537 -1333 -6533
rect -1323 -6537 -1319 -6533
rect -768 -6536 -763 -6532
rect -754 -6536 -750 -6532
rect -745 -6536 -740 -6532
rect -731 -6536 -727 -6532
rect -714 -6536 -710 -6532
rect -700 -6536 -696 -6532
rect -691 -6536 -687 -6532
rect -677 -6536 -673 -6532
rect -613 -6535 -608 -6531
rect -599 -6535 -595 -6531
rect -590 -6535 -585 -6531
rect -576 -6535 -572 -6531
rect -559 -6535 -555 -6531
rect -545 -6535 -541 -6531
rect -536 -6535 -532 -6531
rect -522 -6535 -518 -6531
rect 135 -6536 140 -6532
rect 149 -6536 153 -6532
rect 158 -6536 163 -6532
rect 172 -6536 176 -6532
rect 189 -6536 193 -6532
rect 203 -6536 207 -6532
rect 212 -6536 216 -6532
rect 226 -6536 230 -6532
rect 290 -6535 295 -6531
rect 304 -6535 308 -6531
rect 313 -6535 318 -6531
rect 327 -6535 331 -6531
rect 344 -6535 348 -6531
rect 358 -6535 362 -6531
rect 367 -6535 371 -6531
rect 381 -6535 385 -6531
rect 1003 -6535 1008 -6531
rect 1017 -6535 1021 -6531
rect 1026 -6535 1031 -6531
rect 1040 -6535 1044 -6531
rect 1057 -6535 1061 -6531
rect 1071 -6535 1075 -6531
rect 1080 -6535 1084 -6531
rect 1094 -6535 1098 -6531
rect 1158 -6534 1163 -6530
rect 1172 -6534 1176 -6530
rect 1181 -6534 1186 -6530
rect 1195 -6534 1199 -6530
rect 1212 -6534 1216 -6530
rect 1226 -6534 1230 -6530
rect 1235 -6534 1239 -6530
rect 1249 -6534 1253 -6530
rect 2083 -6510 2088 -6506
rect 2097 -6510 2101 -6506
rect 2106 -6510 2111 -6506
rect 2120 -6510 2124 -6506
rect 2137 -6510 2141 -6506
rect 2151 -6510 2155 -6506
rect 2160 -6510 2164 -6506
rect 2174 -6510 2178 -6506
rect 2217 -6488 2221 -6483
rect 2231 -6488 2235 -6483
rect -1229 -6665 -1225 -6660
rect -1215 -6665 -1211 -6660
rect -1206 -6665 -1202 -6660
rect -1192 -6665 -1188 -6660
rect -1183 -6665 -1179 -6660
rect -1169 -6665 -1165 -6660
rect -1160 -6665 -1156 -6660
rect -1146 -6665 -1142 -6660
rect -428 -6663 -424 -6658
rect -414 -6663 -410 -6658
rect -405 -6663 -401 -6658
rect -391 -6663 -387 -6658
rect -382 -6663 -378 -6658
rect -368 -6663 -364 -6658
rect -359 -6663 -355 -6658
rect -345 -6663 -341 -6658
rect -1675 -6672 -1671 -6667
rect -1661 -6672 -1657 -6667
rect -1652 -6672 -1648 -6667
rect -1638 -6672 -1634 -6667
rect -1614 -6672 -1610 -6667
rect -1600 -6672 -1596 -6667
rect -1535 -6671 -1531 -6666
rect -1521 -6671 -1517 -6666
rect -1512 -6671 -1508 -6666
rect -1498 -6671 -1494 -6666
rect -1474 -6671 -1470 -6666
rect -1460 -6671 -1456 -6666
rect -1390 -6670 -1386 -6665
rect -1376 -6670 -1372 -6665
rect -1367 -6670 -1363 -6665
rect -1353 -6670 -1349 -6665
rect -1329 -6670 -1325 -6665
rect -1315 -6670 -1311 -6665
rect -874 -6670 -870 -6665
rect -860 -6670 -856 -6665
rect -851 -6670 -847 -6665
rect -837 -6670 -833 -6665
rect -813 -6670 -809 -6665
rect -799 -6670 -795 -6665
rect -734 -6669 -730 -6664
rect -720 -6669 -716 -6664
rect -711 -6669 -707 -6664
rect -697 -6669 -693 -6664
rect -673 -6669 -669 -6664
rect -659 -6669 -655 -6664
rect -589 -6668 -585 -6663
rect -575 -6668 -571 -6663
rect -566 -6668 -562 -6663
rect -552 -6668 -548 -6663
rect -528 -6668 -524 -6663
rect -514 -6668 -510 -6663
rect 475 -6663 479 -6658
rect 489 -6663 493 -6658
rect 498 -6663 502 -6658
rect 512 -6663 516 -6658
rect 521 -6663 525 -6658
rect 535 -6663 539 -6658
rect 544 -6663 548 -6658
rect 558 -6663 562 -6658
rect 29 -6670 33 -6665
rect 43 -6670 47 -6665
rect 52 -6670 56 -6665
rect 66 -6670 70 -6665
rect 90 -6670 94 -6665
rect 104 -6670 108 -6665
rect 169 -6669 173 -6664
rect 183 -6669 187 -6664
rect 192 -6669 196 -6664
rect 206 -6669 210 -6664
rect 230 -6669 234 -6664
rect 244 -6669 248 -6664
rect 314 -6668 318 -6663
rect 328 -6668 332 -6663
rect 337 -6668 341 -6663
rect 351 -6668 355 -6663
rect 375 -6668 379 -6663
rect 389 -6668 393 -6663
rect 1343 -6662 1347 -6657
rect 1357 -6662 1361 -6657
rect 1366 -6662 1370 -6657
rect 1380 -6662 1384 -6657
rect 1389 -6662 1393 -6657
rect 1403 -6662 1407 -6657
rect 1412 -6662 1416 -6657
rect 1426 -6662 1430 -6657
rect 897 -6669 901 -6664
rect 911 -6669 915 -6664
rect 920 -6669 924 -6664
rect 934 -6669 938 -6664
rect 958 -6669 962 -6664
rect 972 -6669 976 -6664
rect 1037 -6668 1041 -6663
rect 1051 -6668 1055 -6663
rect 1060 -6668 1064 -6663
rect 1074 -6668 1078 -6663
rect 1098 -6668 1102 -6663
rect 1112 -6668 1116 -6663
rect 1182 -6667 1186 -6662
rect 1196 -6667 1200 -6662
rect 1205 -6667 1209 -6662
rect 1219 -6667 1223 -6662
rect 1243 -6667 1247 -6662
rect 1257 -6667 1261 -6662
rect 3099 -6682 3103 -6677
rect 3113 -6682 3117 -6677
rect 3122 -6682 3126 -6677
rect 3136 -6682 3140 -6677
rect 3145 -6682 3149 -6677
rect 3159 -6682 3163 -6677
rect 3168 -6682 3172 -6677
rect 3182 -6682 3186 -6677
rect 3191 -6682 3195 -6677
rect 3205 -6682 3209 -6677
rect 2088 -6698 2092 -6693
rect 2102 -6698 2106 -6693
rect 2135 -6697 2139 -6692
rect 2149 -6697 2153 -6692
rect 2158 -6697 2162 -6692
rect 2172 -6697 2176 -6692
rect 2214 -6697 2218 -6692
rect 2228 -6697 2232 -6692
rect 2279 -6697 2283 -6692
rect 2293 -6697 2297 -6692
rect 2344 -6697 2348 -6692
rect 2358 -6697 2362 -6692
rect 2367 -6697 2371 -6692
rect 2381 -6697 2385 -6692
rect 2390 -6697 2394 -6692
rect 2404 -6697 2408 -6692
rect 2446 -6697 2450 -6692
rect 2460 -6697 2464 -6692
rect 2506 -6697 2510 -6692
rect 2520 -6697 2524 -6692
rect 2590 -6697 2594 -6692
rect 2604 -6697 2608 -6692
rect 2613 -6697 2617 -6692
rect 2627 -6697 2631 -6692
rect 2636 -6697 2640 -6692
rect 2650 -6697 2654 -6692
rect 2659 -6697 2663 -6692
rect 2673 -6697 2677 -6692
rect 2715 -6697 2719 -6692
rect 2729 -6697 2733 -6692
rect 2777 -6697 2781 -6692
rect 2791 -6697 2795 -6692
rect 2867 -6696 2871 -6691
rect 2881 -6696 2885 -6691
rect 2890 -6696 2894 -6691
rect 2904 -6696 2908 -6691
rect 2913 -6696 2917 -6691
rect 2927 -6696 2931 -6691
rect 2936 -6696 2940 -6691
rect 2950 -6696 2954 -6691
rect 2959 -6696 2963 -6691
rect 2973 -6696 2977 -6691
rect 3015 -6696 3019 -6691
rect 3029 -6696 3033 -6691
<< pdcontact >>
rect 661 -5016 666 -5010
rect 675 -5016 679 -5010
rect 684 -5016 689 -5010
rect 698 -5016 702 -5010
rect 722 -5016 727 -5010
rect 736 -5016 740 -5010
rect 1113 -5101 1118 -5095
rect 1127 -5101 1131 -5095
rect 965 -5118 970 -5112
rect 979 -5118 983 -5112
rect 988 -5118 993 -5112
rect 1002 -5118 1006 -5112
rect 1026 -5118 1031 -5112
rect 1040 -5118 1044 -5112
rect 1203 -5114 1208 -5108
rect 1217 -5114 1221 -5108
rect 1226 -5114 1231 -5108
rect 1240 -5114 1244 -5108
rect 1264 -5114 1269 -5108
rect 1278 -5114 1282 -5108
rect 1334 -5114 1339 -5108
rect 1348 -5114 1352 -5108
rect 1357 -5114 1362 -5108
rect 1371 -5114 1375 -5108
rect 1395 -5114 1400 -5108
rect 1409 -5114 1413 -5108
rect 1490 -5114 1495 -5108
rect 1504 -5114 1508 -5108
rect 1513 -5114 1518 -5108
rect 1527 -5114 1531 -5108
rect 1551 -5114 1556 -5108
rect 1565 -5114 1569 -5108
rect 1112 -5169 1117 -5163
rect 1126 -5169 1130 -5163
rect 567 -5326 572 -5320
rect 581 -5326 585 -5320
rect 590 -5326 595 -5320
rect 604 -5326 608 -5320
rect 633 -5326 638 -5320
rect 647 -5326 651 -5320
rect 675 -5326 680 -5320
rect 689 -5326 693 -5320
rect 698 -5326 703 -5320
rect 712 -5326 716 -5320
rect 741 -5326 746 -5320
rect 755 -5326 759 -5320
rect 787 -5326 792 -5320
rect 801 -5326 805 -5320
rect 810 -5326 815 -5320
rect 824 -5326 828 -5320
rect 853 -5326 858 -5320
rect 867 -5326 871 -5320
rect 899 -5326 904 -5320
rect 913 -5326 917 -5320
rect 922 -5326 927 -5320
rect 936 -5326 940 -5320
rect 965 -5326 970 -5320
rect 979 -5326 983 -5320
rect 1010 -5326 1015 -5320
rect 1024 -5326 1028 -5320
rect 1033 -5326 1038 -5320
rect 1047 -5326 1051 -5320
rect 1076 -5326 1081 -5320
rect 1090 -5326 1094 -5320
rect 1122 -5326 1127 -5320
rect 1136 -5326 1140 -5320
rect 1145 -5326 1150 -5320
rect 1159 -5326 1163 -5320
rect 1188 -5326 1193 -5320
rect 1202 -5326 1206 -5320
rect 1234 -5326 1239 -5320
rect 1248 -5326 1252 -5320
rect 1257 -5326 1262 -5320
rect 1271 -5326 1275 -5320
rect 1300 -5326 1305 -5320
rect 1314 -5326 1318 -5320
rect 1346 -5326 1351 -5320
rect 1360 -5326 1364 -5320
rect 1369 -5326 1374 -5320
rect 1383 -5326 1387 -5320
rect 1412 -5326 1417 -5320
rect 1426 -5326 1430 -5320
rect 1786 -5324 1791 -5318
rect 1800 -5324 1804 -5318
rect 1809 -5324 1814 -5318
rect 1823 -5324 1827 -5318
rect 1852 -5324 1857 -5318
rect 1866 -5324 1870 -5318
rect 1894 -5324 1899 -5318
rect 1908 -5324 1912 -5318
rect 1917 -5324 1922 -5318
rect 1931 -5324 1935 -5318
rect 1960 -5324 1965 -5318
rect 1974 -5324 1978 -5318
rect 2006 -5324 2011 -5318
rect 2020 -5324 2024 -5318
rect 2029 -5324 2034 -5318
rect 2043 -5324 2047 -5318
rect 2072 -5324 2077 -5318
rect 2086 -5324 2090 -5318
rect 2118 -5324 2123 -5318
rect 2132 -5324 2136 -5318
rect 2141 -5324 2146 -5318
rect 2155 -5324 2159 -5318
rect 2184 -5324 2189 -5318
rect 2198 -5324 2202 -5318
rect 2229 -5324 2234 -5318
rect 2243 -5324 2247 -5318
rect 2252 -5324 2257 -5318
rect 2266 -5324 2270 -5318
rect 2295 -5324 2300 -5318
rect 2309 -5324 2313 -5318
rect 2341 -5324 2346 -5318
rect 2355 -5324 2359 -5318
rect 2364 -5324 2369 -5318
rect 2378 -5324 2382 -5318
rect 2407 -5324 2412 -5318
rect 2421 -5324 2425 -5318
rect 2453 -5324 2458 -5318
rect 2467 -5324 2471 -5318
rect 2476 -5324 2481 -5318
rect 2490 -5324 2494 -5318
rect 2519 -5324 2524 -5318
rect 2533 -5324 2537 -5318
rect 2565 -5324 2570 -5318
rect 2579 -5324 2583 -5318
rect 2588 -5324 2593 -5318
rect 2602 -5324 2606 -5318
rect 2631 -5324 2636 -5318
rect 2645 -5324 2649 -5318
rect -584 -5333 -579 -5327
rect -570 -5333 -566 -5327
rect -561 -5333 -556 -5327
rect -547 -5333 -543 -5327
rect -518 -5333 -513 -5327
rect -504 -5333 -500 -5327
rect -476 -5333 -471 -5327
rect -462 -5333 -458 -5327
rect -453 -5333 -448 -5327
rect -439 -5333 -435 -5327
rect -410 -5333 -405 -5327
rect -396 -5333 -392 -5327
rect -364 -5333 -359 -5327
rect -350 -5333 -346 -5327
rect -341 -5333 -336 -5327
rect -327 -5333 -323 -5327
rect -298 -5333 -293 -5327
rect -284 -5333 -280 -5327
rect -252 -5333 -247 -5327
rect -238 -5333 -234 -5327
rect -229 -5333 -224 -5327
rect -215 -5333 -211 -5327
rect -186 -5333 -181 -5327
rect -172 -5333 -168 -5327
rect -141 -5333 -136 -5327
rect -127 -5333 -123 -5327
rect -118 -5333 -113 -5327
rect -104 -5333 -100 -5327
rect -75 -5333 -70 -5327
rect -61 -5333 -57 -5327
rect -29 -5333 -24 -5327
rect -15 -5333 -11 -5327
rect -6 -5333 -1 -5327
rect 8 -5333 12 -5327
rect 37 -5333 42 -5327
rect 51 -5333 55 -5327
rect 83 -5333 88 -5327
rect 97 -5333 101 -5327
rect 106 -5333 111 -5327
rect 120 -5333 124 -5327
rect 149 -5333 154 -5327
rect 163 -5333 167 -5327
rect 195 -5333 200 -5327
rect 209 -5333 213 -5327
rect 218 -5333 223 -5327
rect 232 -5333 236 -5327
rect 261 -5333 266 -5327
rect 275 -5333 279 -5327
rect 2569 -5715 2574 -5709
rect 2583 -5715 2587 -5709
rect 2592 -5715 2597 -5709
rect 2606 -5715 2610 -5709
rect 2615 -5715 2620 -5709
rect 2629 -5715 2633 -5709
rect 2638 -5715 2643 -5709
rect 2652 -5715 2656 -5709
rect 2661 -5715 2666 -5709
rect 2675 -5715 2679 -5709
rect -550 -5817 -545 -5811
rect -536 -5817 -532 -5811
rect -527 -5817 -522 -5811
rect -513 -5817 -509 -5811
rect -489 -5817 -484 -5811
rect -475 -5817 -471 -5811
rect -411 -5817 -406 -5811
rect -397 -5817 -393 -5811
rect -388 -5817 -383 -5811
rect -374 -5817 -370 -5811
rect -350 -5817 -345 -5811
rect -336 -5817 -332 -5811
rect -273 -5817 -268 -5811
rect -259 -5817 -255 -5811
rect -250 -5817 -245 -5811
rect -236 -5817 -232 -5811
rect -212 -5817 -207 -5811
rect -198 -5817 -194 -5811
rect -123 -5817 -118 -5811
rect -109 -5817 -105 -5811
rect -100 -5817 -95 -5811
rect -86 -5817 -82 -5811
rect -62 -5817 -57 -5811
rect -48 -5817 -44 -5811
rect 2141 -5853 2146 -5847
rect 2155 -5853 2159 -5847
rect 2164 -5853 2169 -5847
rect 2178 -5853 2182 -5847
rect 2220 -5853 2225 -5847
rect 2234 -5853 2238 -5847
rect 2342 -5853 2347 -5847
rect 2356 -5853 2360 -5847
rect 2365 -5853 2370 -5847
rect 2379 -5853 2383 -5847
rect 2388 -5853 2393 -5847
rect 2402 -5853 2406 -5847
rect 2444 -5853 2449 -5847
rect 2458 -5853 2462 -5847
rect 2589 -5853 2594 -5847
rect 2603 -5853 2607 -5847
rect 2612 -5853 2617 -5847
rect 2626 -5853 2630 -5847
rect 2635 -5853 2640 -5847
rect 2649 -5853 2653 -5847
rect 2658 -5853 2663 -5847
rect 2672 -5853 2676 -5847
rect 2714 -5853 2719 -5847
rect 2728 -5853 2732 -5847
rect 2869 -5853 2874 -5847
rect 2883 -5853 2887 -5847
rect 2892 -5853 2897 -5847
rect 2906 -5853 2910 -5847
rect 2915 -5853 2920 -5847
rect 2929 -5853 2933 -5847
rect 2938 -5853 2943 -5847
rect 2952 -5853 2956 -5847
rect 2961 -5853 2966 -5847
rect 2975 -5853 2979 -5847
rect 3017 -5853 3022 -5847
rect 3031 -5853 3035 -5847
rect 2094 -5864 2099 -5858
rect 2108 -5864 2112 -5858
rect 2277 -5863 2282 -5857
rect 2291 -5863 2295 -5857
rect 2505 -5863 2510 -5857
rect 2519 -5863 2523 -5857
rect 2779 -5864 2784 -5858
rect 2793 -5864 2797 -5858
rect 2083 -5996 2088 -5990
rect 2097 -5996 2101 -5990
rect 2106 -5996 2111 -5990
rect 2120 -5996 2124 -5990
rect 2137 -5996 2142 -5990
rect 2151 -5996 2155 -5990
rect 2160 -5996 2165 -5990
rect 2174 -5996 2178 -5990
rect 2217 -6001 2222 -5995
rect 2231 -6001 2235 -5995
rect -1582 -6174 -1577 -6168
rect -1568 -6174 -1564 -6168
rect -1559 -6174 -1554 -6168
rect -1545 -6174 -1541 -6168
rect -1528 -6174 -1523 -6168
rect -1514 -6174 -1510 -6168
rect -1505 -6174 -1500 -6168
rect -1491 -6174 -1487 -6168
rect -792 -6174 -787 -6168
rect -778 -6174 -774 -6168
rect -769 -6174 -764 -6168
rect -755 -6174 -751 -6168
rect -738 -6174 -733 -6168
rect -724 -6174 -720 -6168
rect -715 -6174 -710 -6168
rect -701 -6174 -697 -6168
rect 190 -6174 195 -6168
rect 204 -6174 208 -6168
rect 213 -6174 218 -6168
rect 227 -6174 231 -6168
rect 244 -6174 249 -6168
rect 258 -6174 262 -6168
rect 267 -6174 272 -6168
rect 281 -6174 285 -6168
rect 1074 -6174 1079 -6168
rect 1088 -6174 1092 -6168
rect 1097 -6174 1102 -6168
rect 1111 -6174 1115 -6168
rect 1128 -6174 1133 -6168
rect 1142 -6174 1146 -6168
rect 1151 -6174 1156 -6168
rect 1165 -6174 1169 -6168
rect 2082 -6141 2087 -6135
rect 2096 -6141 2100 -6135
rect 2105 -6141 2110 -6135
rect 2119 -6141 2123 -6135
rect 2136 -6141 2141 -6135
rect 2150 -6141 2154 -6135
rect 2159 -6141 2164 -6135
rect 2173 -6141 2177 -6135
rect 2216 -6146 2221 -6140
rect 2230 -6146 2234 -6140
rect 2346 -6228 2351 -6222
rect 2360 -6228 2364 -6222
rect 2369 -6228 2374 -6222
rect 2383 -6228 2387 -6222
rect 2392 -6228 2397 -6222
rect 2406 -6228 2410 -6222
rect 2415 -6228 2420 -6222
rect 2429 -6228 2433 -6222
rect 2471 -6228 2476 -6222
rect 2485 -6228 2489 -6222
rect 2082 -6303 2087 -6297
rect 2096 -6303 2100 -6297
rect 2105 -6303 2110 -6297
rect 2119 -6303 2123 -6297
rect 2136 -6303 2141 -6297
rect 2150 -6303 2154 -6297
rect 2159 -6303 2164 -6297
rect 2173 -6303 2177 -6297
rect 2216 -6308 2221 -6302
rect 2230 -6308 2234 -6302
rect -1569 -6485 -1564 -6479
rect -1555 -6485 -1551 -6479
rect -1546 -6485 -1541 -6479
rect -1532 -6485 -1528 -6479
rect -1515 -6485 -1510 -6479
rect -1501 -6485 -1497 -6479
rect -1492 -6485 -1487 -6479
rect -1478 -6485 -1474 -6479
rect -1414 -6484 -1409 -6478
rect -1400 -6484 -1396 -6478
rect -1391 -6484 -1386 -6478
rect -1377 -6484 -1373 -6478
rect -1360 -6484 -1355 -6478
rect -1346 -6484 -1342 -6478
rect -1337 -6484 -1332 -6478
rect -1323 -6484 -1319 -6478
rect -768 -6483 -763 -6477
rect -754 -6483 -750 -6477
rect -745 -6483 -740 -6477
rect -731 -6483 -727 -6477
rect -714 -6483 -709 -6477
rect -700 -6483 -696 -6477
rect -691 -6483 -686 -6477
rect -677 -6483 -673 -6477
rect -613 -6482 -608 -6476
rect -599 -6482 -595 -6476
rect -590 -6482 -585 -6476
rect -576 -6482 -572 -6476
rect -559 -6482 -554 -6476
rect -545 -6482 -541 -6476
rect -536 -6482 -531 -6476
rect -522 -6482 -518 -6476
rect 135 -6483 140 -6477
rect 149 -6483 153 -6477
rect 158 -6483 163 -6477
rect 172 -6483 176 -6477
rect 189 -6483 194 -6477
rect 203 -6483 207 -6477
rect 212 -6483 217 -6477
rect 226 -6483 230 -6477
rect 290 -6482 295 -6476
rect 304 -6482 308 -6476
rect 313 -6482 318 -6476
rect 327 -6482 331 -6476
rect 344 -6482 349 -6476
rect 358 -6482 362 -6476
rect 367 -6482 372 -6476
rect 381 -6482 385 -6476
rect 1003 -6482 1008 -6476
rect 1017 -6482 1021 -6476
rect 1026 -6482 1031 -6476
rect 1040 -6482 1044 -6476
rect 1057 -6482 1062 -6476
rect 1071 -6482 1075 -6476
rect 1080 -6482 1085 -6476
rect 1094 -6482 1098 -6476
rect 1158 -6481 1163 -6475
rect 1172 -6481 1176 -6475
rect 1181 -6481 1186 -6475
rect 1195 -6481 1199 -6475
rect 1212 -6481 1217 -6475
rect 1226 -6481 1230 -6475
rect 1235 -6481 1240 -6475
rect 1249 -6481 1253 -6475
rect 2083 -6457 2088 -6451
rect 2097 -6457 2101 -6451
rect 2106 -6457 2111 -6451
rect 2120 -6457 2124 -6451
rect 2137 -6457 2142 -6451
rect 2151 -6457 2155 -6451
rect 2160 -6457 2165 -6451
rect 2174 -6457 2178 -6451
rect 2217 -6462 2222 -6456
rect 2231 -6462 2235 -6456
rect -1675 -6636 -1670 -6630
rect -1661 -6636 -1657 -6630
rect -1652 -6636 -1647 -6630
rect -1638 -6636 -1634 -6630
rect -1614 -6636 -1609 -6630
rect -1600 -6636 -1596 -6630
rect -1535 -6635 -1530 -6629
rect -1521 -6635 -1517 -6629
rect -1512 -6635 -1507 -6629
rect -1498 -6635 -1494 -6629
rect -1474 -6635 -1469 -6629
rect -1460 -6635 -1456 -6629
rect -1390 -6634 -1385 -6628
rect -1376 -6634 -1372 -6628
rect -1367 -6634 -1362 -6628
rect -1353 -6634 -1349 -6628
rect -1329 -6634 -1324 -6628
rect -1315 -6634 -1311 -6628
rect -1229 -6637 -1224 -6631
rect -1215 -6637 -1211 -6631
rect -1206 -6637 -1201 -6631
rect -1192 -6637 -1188 -6631
rect -1183 -6637 -1178 -6631
rect -1169 -6637 -1165 -6631
rect -1160 -6637 -1155 -6631
rect -1146 -6637 -1142 -6631
rect -874 -6634 -869 -6628
rect -860 -6634 -856 -6628
rect -851 -6634 -846 -6628
rect -837 -6634 -833 -6628
rect -813 -6634 -808 -6628
rect -799 -6634 -795 -6628
rect -734 -6633 -729 -6627
rect -720 -6633 -716 -6627
rect -711 -6633 -706 -6627
rect -697 -6633 -693 -6627
rect -673 -6633 -668 -6627
rect -659 -6633 -655 -6627
rect -589 -6632 -584 -6626
rect -575 -6632 -571 -6626
rect -566 -6632 -561 -6626
rect -552 -6632 -548 -6626
rect -528 -6632 -523 -6626
rect -514 -6632 -510 -6626
rect -428 -6635 -423 -6629
rect -414 -6635 -410 -6629
rect -405 -6635 -400 -6629
rect -391 -6635 -387 -6629
rect -382 -6635 -377 -6629
rect -368 -6635 -364 -6629
rect -359 -6635 -354 -6629
rect -345 -6635 -341 -6629
rect 29 -6634 34 -6628
rect 43 -6634 47 -6628
rect 52 -6634 57 -6628
rect 66 -6634 70 -6628
rect 90 -6634 95 -6628
rect 104 -6634 108 -6628
rect 169 -6633 174 -6627
rect 183 -6633 187 -6627
rect 192 -6633 197 -6627
rect 206 -6633 210 -6627
rect 230 -6633 235 -6627
rect 244 -6633 248 -6627
rect 314 -6632 319 -6626
rect 328 -6632 332 -6626
rect 337 -6632 342 -6626
rect 351 -6632 355 -6626
rect 375 -6632 380 -6626
rect 389 -6632 393 -6626
rect 475 -6635 480 -6629
rect 489 -6635 493 -6629
rect 498 -6635 503 -6629
rect 512 -6635 516 -6629
rect 521 -6635 526 -6629
rect 535 -6635 539 -6629
rect 544 -6635 549 -6629
rect 558 -6635 562 -6629
rect 897 -6633 902 -6627
rect 911 -6633 915 -6627
rect 920 -6633 925 -6627
rect 934 -6633 938 -6627
rect 958 -6633 963 -6627
rect 972 -6633 976 -6627
rect 1037 -6632 1042 -6626
rect 1051 -6632 1055 -6626
rect 1060 -6632 1065 -6626
rect 1074 -6632 1078 -6626
rect 1098 -6632 1103 -6626
rect 1112 -6632 1116 -6626
rect 1182 -6631 1187 -6625
rect 1196 -6631 1200 -6625
rect 1205 -6631 1210 -6625
rect 1219 -6631 1223 -6625
rect 1243 -6631 1248 -6625
rect 1257 -6631 1261 -6625
rect 1343 -6634 1348 -6628
rect 1357 -6634 1361 -6628
rect 1366 -6634 1371 -6628
rect 1380 -6634 1384 -6628
rect 1389 -6634 1394 -6628
rect 1403 -6634 1407 -6628
rect 1412 -6634 1417 -6628
rect 1426 -6634 1430 -6628
rect 3099 -6654 3104 -6648
rect 3113 -6654 3117 -6648
rect 3122 -6654 3127 -6648
rect 3136 -6654 3140 -6648
rect 3145 -6654 3150 -6648
rect 3159 -6654 3163 -6648
rect 3168 -6654 3173 -6648
rect 3182 -6654 3186 -6648
rect 3191 -6654 3196 -6648
rect 3205 -6654 3209 -6648
rect 2135 -6661 2140 -6655
rect 2149 -6661 2153 -6655
rect 2158 -6661 2163 -6655
rect 2172 -6661 2176 -6655
rect 2214 -6661 2219 -6655
rect 2228 -6661 2232 -6655
rect 2344 -6661 2349 -6655
rect 2358 -6661 2362 -6655
rect 2367 -6661 2372 -6655
rect 2381 -6661 2385 -6655
rect 2390 -6661 2395 -6655
rect 2404 -6661 2408 -6655
rect 2446 -6661 2451 -6655
rect 2460 -6661 2464 -6655
rect 2590 -6661 2595 -6655
rect 2604 -6661 2608 -6655
rect 2613 -6661 2618 -6655
rect 2627 -6661 2631 -6655
rect 2636 -6661 2641 -6655
rect 2650 -6661 2654 -6655
rect 2659 -6661 2664 -6655
rect 2673 -6661 2677 -6655
rect 2715 -6661 2720 -6655
rect 2729 -6661 2733 -6655
rect 2867 -6660 2872 -6654
rect 2881 -6660 2885 -6654
rect 2890 -6660 2895 -6654
rect 2904 -6660 2908 -6654
rect 2913 -6660 2918 -6654
rect 2927 -6660 2931 -6654
rect 2936 -6660 2941 -6654
rect 2950 -6660 2954 -6654
rect 2959 -6660 2964 -6654
rect 2973 -6660 2977 -6654
rect 3015 -6660 3020 -6654
rect 3029 -6660 3033 -6654
rect 2088 -6672 2093 -6666
rect 2102 -6672 2106 -6666
rect 2279 -6671 2284 -6665
rect 2293 -6671 2297 -6665
rect 2506 -6671 2511 -6665
rect 2520 -6671 2524 -6665
rect 2777 -6671 2782 -6665
rect 2791 -6671 2795 -6665
<< polysilicon >>
rect 669 -5010 672 -5007
rect 692 -5010 695 -5007
rect 730 -5010 733 -5007
rect 669 -5047 672 -5016
rect 692 -5037 695 -5016
rect 730 -5026 733 -5016
rect 728 -5030 733 -5026
rect 690 -5041 695 -5037
rect 692 -5047 695 -5041
rect 730 -5047 733 -5030
rect 669 -5056 672 -5052
rect 692 -5056 695 -5052
rect 730 -5056 733 -5052
rect 1121 -5095 1124 -5092
rect 973 -5112 976 -5109
rect 996 -5112 999 -5109
rect 1034 -5112 1037 -5109
rect 1121 -5112 1124 -5101
rect 1211 -5108 1214 -5105
rect 1234 -5108 1237 -5105
rect 1272 -5108 1275 -5105
rect 1342 -5108 1345 -5105
rect 1365 -5108 1368 -5105
rect 1403 -5108 1406 -5105
rect 1498 -5108 1501 -5105
rect 1521 -5108 1524 -5105
rect 1559 -5108 1562 -5105
rect 1119 -5116 1124 -5112
rect 973 -5149 976 -5118
rect 996 -5139 999 -5118
rect 1034 -5128 1037 -5118
rect 1121 -5122 1124 -5116
rect 1211 -5125 1214 -5114
rect 1032 -5132 1037 -5128
rect 994 -5143 999 -5139
rect 996 -5149 999 -5143
rect 1034 -5149 1037 -5132
rect 1121 -5134 1124 -5127
rect 1209 -5129 1214 -5125
rect 1211 -5145 1214 -5129
rect 1234 -5134 1237 -5114
rect 1272 -5124 1275 -5114
rect 1270 -5128 1275 -5124
rect 1342 -5125 1345 -5114
rect 1232 -5138 1237 -5134
rect 1234 -5145 1237 -5138
rect 1272 -5145 1275 -5128
rect 1340 -5129 1345 -5125
rect 1342 -5145 1345 -5129
rect 1365 -5134 1368 -5114
rect 1403 -5124 1406 -5114
rect 1401 -5128 1406 -5124
rect 1498 -5125 1501 -5114
rect 1363 -5138 1368 -5134
rect 1365 -5145 1368 -5138
rect 1403 -5145 1406 -5128
rect 1496 -5129 1501 -5125
rect 1498 -5145 1501 -5129
rect 1521 -5134 1524 -5114
rect 1559 -5124 1562 -5114
rect 1557 -5128 1562 -5124
rect 1519 -5138 1524 -5134
rect 1521 -5145 1524 -5138
rect 1559 -5145 1562 -5128
rect 1211 -5154 1214 -5150
rect 1234 -5154 1237 -5150
rect 1272 -5154 1275 -5150
rect 1342 -5154 1345 -5150
rect 1365 -5154 1368 -5150
rect 1403 -5154 1406 -5150
rect 1498 -5154 1501 -5150
rect 1521 -5154 1524 -5150
rect 1559 -5154 1562 -5150
rect 973 -5158 976 -5154
rect 996 -5158 999 -5154
rect 1034 -5158 1037 -5154
rect 1120 -5163 1123 -5160
rect 1120 -5180 1123 -5169
rect 1118 -5184 1123 -5180
rect 1120 -5190 1123 -5184
rect 1120 -5202 1123 -5195
rect -576 -5327 -573 -5308
rect -553 -5327 -550 -5324
rect -510 -5327 -507 -5324
rect -468 -5327 -465 -5308
rect -445 -5327 -442 -5324
rect -402 -5327 -399 -5324
rect -356 -5327 -353 -5308
rect -333 -5327 -330 -5324
rect -290 -5327 -287 -5324
rect -244 -5327 -241 -5308
rect -221 -5327 -218 -5324
rect -178 -5327 -175 -5324
rect -133 -5327 -130 -5308
rect -110 -5327 -107 -5324
rect -67 -5327 -64 -5324
rect -21 -5327 -18 -5308
rect 2 -5327 5 -5324
rect 45 -5327 48 -5324
rect 91 -5327 94 -5308
rect 114 -5327 117 -5324
rect 157 -5327 160 -5324
rect 203 -5327 206 -5308
rect 575 -5320 578 -5301
rect 598 -5320 601 -5317
rect 641 -5320 644 -5317
rect 683 -5320 686 -5301
rect 706 -5320 709 -5317
rect 749 -5320 752 -5317
rect 795 -5320 798 -5301
rect 818 -5320 821 -5317
rect 861 -5320 864 -5317
rect 907 -5320 910 -5301
rect 930 -5320 933 -5317
rect 973 -5320 976 -5317
rect 1018 -5320 1021 -5301
rect 1041 -5320 1044 -5317
rect 1084 -5320 1087 -5317
rect 1130 -5320 1133 -5301
rect 1153 -5320 1156 -5317
rect 1196 -5320 1199 -5317
rect 1242 -5320 1245 -5301
rect 1265 -5320 1268 -5317
rect 1308 -5320 1311 -5317
rect 1354 -5320 1357 -5301
rect 1377 -5320 1380 -5317
rect 1420 -5320 1423 -5317
rect 1794 -5318 1797 -5299
rect 1817 -5318 1820 -5315
rect 1860 -5318 1863 -5315
rect 1902 -5318 1905 -5299
rect 1925 -5318 1928 -5315
rect 1968 -5318 1971 -5315
rect 2014 -5318 2017 -5299
rect 2037 -5318 2040 -5315
rect 2080 -5318 2083 -5315
rect 2126 -5318 2129 -5299
rect 2149 -5318 2152 -5315
rect 2192 -5318 2195 -5315
rect 2237 -5318 2240 -5299
rect 2260 -5318 2263 -5315
rect 2303 -5318 2306 -5315
rect 2349 -5318 2352 -5299
rect 2372 -5318 2375 -5315
rect 2415 -5318 2418 -5315
rect 2461 -5318 2464 -5299
rect 2484 -5318 2487 -5315
rect 2527 -5318 2530 -5315
rect 2573 -5318 2576 -5299
rect 2596 -5318 2599 -5315
rect 2639 -5318 2642 -5315
rect 226 -5327 229 -5324
rect 269 -5327 272 -5324
rect -576 -5364 -573 -5333
rect -553 -5364 -550 -5333
rect -510 -5343 -507 -5333
rect -512 -5347 -507 -5343
rect -510 -5364 -507 -5347
rect -468 -5364 -465 -5333
rect -445 -5364 -442 -5333
rect -402 -5343 -399 -5333
rect -404 -5347 -399 -5343
rect -402 -5364 -399 -5347
rect -356 -5364 -353 -5333
rect -333 -5364 -330 -5333
rect -290 -5343 -287 -5333
rect -292 -5347 -287 -5343
rect -290 -5364 -287 -5347
rect -244 -5364 -241 -5333
rect -221 -5364 -218 -5333
rect -178 -5343 -175 -5333
rect -180 -5347 -175 -5343
rect -178 -5364 -175 -5347
rect -133 -5364 -130 -5333
rect -110 -5364 -107 -5333
rect -67 -5343 -64 -5333
rect -69 -5347 -64 -5343
rect -67 -5364 -64 -5347
rect -21 -5364 -18 -5333
rect 2 -5364 5 -5333
rect 45 -5343 48 -5333
rect 43 -5347 48 -5343
rect 45 -5364 48 -5347
rect 91 -5364 94 -5333
rect 114 -5364 117 -5333
rect 157 -5343 160 -5333
rect 155 -5347 160 -5343
rect 157 -5364 160 -5347
rect 203 -5364 206 -5333
rect 226 -5364 229 -5333
rect 269 -5343 272 -5333
rect 267 -5347 272 -5343
rect 269 -5364 272 -5347
rect 575 -5357 578 -5326
rect 598 -5357 601 -5326
rect 641 -5336 644 -5326
rect 639 -5340 644 -5336
rect 641 -5357 644 -5340
rect 683 -5357 686 -5326
rect 706 -5357 709 -5326
rect 749 -5336 752 -5326
rect 747 -5340 752 -5336
rect 749 -5357 752 -5340
rect 795 -5357 798 -5326
rect 818 -5357 821 -5326
rect 861 -5336 864 -5326
rect 859 -5340 864 -5336
rect 861 -5357 864 -5340
rect 907 -5357 910 -5326
rect 930 -5357 933 -5326
rect 973 -5336 976 -5326
rect 971 -5340 976 -5336
rect 973 -5357 976 -5340
rect 1018 -5357 1021 -5326
rect 1041 -5357 1044 -5326
rect 1084 -5336 1087 -5326
rect 1082 -5340 1087 -5336
rect 1084 -5357 1087 -5340
rect 1130 -5357 1133 -5326
rect 1153 -5357 1156 -5326
rect 1196 -5336 1199 -5326
rect 1194 -5340 1199 -5336
rect 1196 -5357 1199 -5340
rect 1242 -5357 1245 -5326
rect 1265 -5357 1268 -5326
rect 1308 -5336 1311 -5326
rect 1306 -5340 1311 -5336
rect 1308 -5357 1311 -5340
rect 1354 -5357 1357 -5326
rect 1377 -5357 1380 -5326
rect 1420 -5336 1423 -5326
rect 1418 -5340 1423 -5336
rect 1420 -5357 1423 -5340
rect 1794 -5355 1797 -5324
rect 1817 -5355 1820 -5324
rect 1860 -5334 1863 -5324
rect 1858 -5338 1863 -5334
rect 1860 -5355 1863 -5338
rect 1902 -5355 1905 -5324
rect 1925 -5355 1928 -5324
rect 1968 -5334 1971 -5324
rect 1966 -5338 1971 -5334
rect 1968 -5355 1971 -5338
rect 2014 -5355 2017 -5324
rect 2037 -5355 2040 -5324
rect 2080 -5334 2083 -5324
rect 2078 -5338 2083 -5334
rect 2080 -5355 2083 -5338
rect 2126 -5355 2129 -5324
rect 2149 -5355 2152 -5324
rect 2192 -5334 2195 -5324
rect 2190 -5338 2195 -5334
rect 2192 -5355 2195 -5338
rect 2237 -5355 2240 -5324
rect 2260 -5355 2263 -5324
rect 2303 -5334 2306 -5324
rect 2301 -5338 2306 -5334
rect 2303 -5355 2306 -5338
rect 2349 -5355 2352 -5324
rect 2372 -5355 2375 -5324
rect 2415 -5334 2418 -5324
rect 2413 -5338 2418 -5334
rect 2415 -5355 2418 -5338
rect 2461 -5355 2464 -5324
rect 2484 -5355 2487 -5324
rect 2527 -5334 2530 -5324
rect 2525 -5338 2530 -5334
rect 2527 -5355 2530 -5338
rect 2573 -5355 2576 -5324
rect 2596 -5355 2599 -5324
rect 2639 -5334 2642 -5324
rect 2637 -5338 2642 -5334
rect 2639 -5355 2642 -5338
rect 575 -5366 578 -5362
rect 598 -5366 601 -5362
rect 641 -5366 644 -5362
rect 683 -5366 686 -5362
rect 706 -5365 709 -5362
rect 581 -5368 601 -5366
rect 695 -5367 709 -5365
rect 749 -5366 752 -5362
rect 795 -5366 798 -5362
rect 818 -5366 821 -5362
rect 861 -5366 864 -5362
rect 907 -5366 910 -5362
rect 930 -5365 933 -5362
rect -576 -5373 -573 -5369
rect -553 -5569 -550 -5369
rect -510 -5374 -507 -5369
rect -468 -5373 -465 -5369
rect -445 -5565 -442 -5369
rect -402 -5373 -399 -5369
rect -356 -5373 -353 -5369
rect -333 -5550 -330 -5369
rect -290 -5373 -287 -5369
rect -244 -5373 -241 -5369
rect -221 -5527 -218 -5369
rect -178 -5373 -175 -5369
rect -133 -5373 -130 -5369
rect -110 -5506 -107 -5369
rect -67 -5373 -64 -5369
rect -21 -5373 -18 -5369
rect 2 -5477 5 -5369
rect 45 -5373 48 -5369
rect 91 -5373 94 -5369
rect 114 -5454 117 -5369
rect 157 -5373 160 -5369
rect 203 -5373 206 -5369
rect 226 -5436 229 -5369
rect 269 -5373 272 -5369
rect -553 -5577 -549 -5569
rect 581 -5579 585 -5368
rect 695 -5377 699 -5367
rect 677 -5380 699 -5377
rect 806 -5368 821 -5366
rect 918 -5367 933 -5365
rect 973 -5366 976 -5362
rect 1018 -5366 1021 -5362
rect 1041 -5366 1044 -5362
rect 1084 -5366 1087 -5362
rect 1130 -5366 1133 -5362
rect 806 -5379 811 -5368
rect 677 -5567 683 -5380
rect 789 -5384 811 -5379
rect 918 -5381 922 -5367
rect 789 -5549 794 -5384
rect 901 -5386 922 -5381
rect 1025 -5368 1044 -5366
rect 1153 -5367 1156 -5362
rect 1196 -5366 1199 -5362
rect 1242 -5366 1245 -5362
rect 1265 -5365 1268 -5362
rect 901 -5525 906 -5386
rect 1025 -5506 1031 -5368
rect 1143 -5369 1156 -5367
rect 1248 -5367 1268 -5365
rect 1308 -5366 1311 -5362
rect 1354 -5366 1357 -5362
rect 1377 -5366 1380 -5362
rect 1420 -5366 1423 -5362
rect 1794 -5364 1797 -5360
rect 1143 -5475 1148 -5369
rect 1248 -5456 1252 -5367
rect 1365 -5368 1380 -5366
rect 1365 -5438 1369 -5368
rect 1143 -5476 1150 -5475
rect 1817 -5569 1820 -5360
rect 1860 -5364 1863 -5360
rect 1902 -5364 1905 -5360
rect 1925 -5566 1928 -5360
rect 1968 -5364 1971 -5360
rect 2014 -5364 2017 -5360
rect 2037 -5364 2040 -5360
rect 2080 -5364 2083 -5360
rect 2126 -5364 2129 -5360
rect 2036 -5551 2040 -5364
rect 2149 -5526 2152 -5360
rect 2192 -5364 2195 -5360
rect 2237 -5364 2240 -5360
rect 2260 -5507 2263 -5360
rect 2303 -5364 2306 -5360
rect 2349 -5364 2352 -5360
rect 2372 -5476 2375 -5360
rect 2415 -5364 2418 -5360
rect 2461 -5364 2464 -5360
rect 2484 -5455 2487 -5360
rect 2527 -5364 2530 -5360
rect 2573 -5364 2576 -5360
rect 2596 -5438 2599 -5360
rect 2639 -5364 2642 -5360
rect 1817 -5578 1821 -5569
rect 2577 -5709 2580 -5705
rect 2600 -5709 2603 -5705
rect 2623 -5709 2626 -5705
rect 2646 -5709 2649 -5705
rect 2669 -5709 2672 -5705
rect 2577 -5738 2580 -5715
rect 2600 -5738 2603 -5715
rect 2623 -5738 2626 -5715
rect 2646 -5738 2649 -5715
rect 2669 -5727 2672 -5715
rect 2667 -5731 2672 -5727
rect 2669 -5738 2672 -5731
rect 2577 -5763 2580 -5743
rect 2600 -5763 2603 -5743
rect 2623 -5763 2626 -5743
rect 2646 -5759 2649 -5743
rect 2669 -5750 2672 -5743
rect -542 -5811 -539 -5789
rect -519 -5811 -516 -5789
rect -481 -5811 -478 -5808
rect -403 -5811 -400 -5788
rect -380 -5811 -377 -5787
rect -342 -5811 -339 -5808
rect -265 -5811 -262 -5788
rect -242 -5811 -239 -5788
rect -204 -5811 -201 -5808
rect -115 -5811 -112 -5787
rect -92 -5811 -89 -5787
rect -54 -5811 -51 -5808
rect -542 -5848 -539 -5817
rect -519 -5848 -516 -5817
rect -481 -5827 -478 -5817
rect -483 -5831 -478 -5827
rect -481 -5848 -478 -5831
rect -403 -5848 -400 -5817
rect -380 -5848 -377 -5817
rect -342 -5827 -339 -5817
rect -344 -5831 -339 -5827
rect -342 -5848 -339 -5831
rect -265 -5848 -262 -5817
rect -242 -5848 -239 -5817
rect -204 -5827 -201 -5817
rect -206 -5831 -201 -5827
rect -204 -5848 -201 -5831
rect -115 -5848 -112 -5817
rect -92 -5848 -89 -5817
rect -54 -5827 -51 -5817
rect -56 -5831 -51 -5827
rect -54 -5848 -51 -5831
rect 2149 -5847 2152 -5844
rect 2172 -5847 2175 -5831
rect 2228 -5847 2231 -5844
rect 2350 -5847 2353 -5844
rect 2373 -5847 2376 -5832
rect 2396 -5847 2399 -5844
rect 2452 -5847 2455 -5844
rect 2597 -5847 2600 -5844
rect 2620 -5847 2623 -5800
rect 2643 -5847 2646 -5844
rect 2666 -5847 2669 -5844
rect 2722 -5847 2725 -5844
rect 2877 -5847 2880 -5844
rect 2900 -5847 2903 -5831
rect 2923 -5847 2926 -5844
rect 2946 -5847 2949 -5844
rect 2969 -5847 2972 -5844
rect 3025 -5847 3028 -5844
rect -542 -5857 -539 -5853
rect -519 -5857 -516 -5853
rect -481 -5857 -478 -5853
rect -403 -5857 -400 -5853
rect -380 -5857 -377 -5853
rect -342 -5857 -339 -5853
rect -265 -5857 -262 -5853
rect -242 -5857 -239 -5853
rect -204 -5857 -201 -5853
rect -115 -5857 -112 -5853
rect -92 -5857 -89 -5853
rect -54 -5857 -51 -5853
rect 2102 -5858 2105 -5855
rect 2102 -5875 2105 -5864
rect 2149 -5873 2152 -5853
rect 2100 -5879 2105 -5875
rect 2147 -5877 2152 -5873
rect 2102 -5885 2105 -5879
rect 2149 -5884 2152 -5877
rect 2172 -5884 2175 -5853
rect 2228 -5863 2231 -5853
rect 2285 -5857 2288 -5854
rect 2350 -5862 2353 -5853
rect 2226 -5867 2231 -5863
rect 2228 -5884 2231 -5867
rect 2285 -5874 2288 -5863
rect 2344 -5866 2353 -5862
rect 2283 -5878 2288 -5874
rect 2285 -5884 2288 -5878
rect 2350 -5884 2353 -5866
rect 2373 -5868 2376 -5853
rect 2371 -5872 2376 -5868
rect 2373 -5884 2376 -5872
rect 2396 -5873 2399 -5853
rect 2452 -5863 2455 -5853
rect 2513 -5857 2516 -5854
rect 2597 -5862 2600 -5853
rect 2450 -5867 2455 -5863
rect 2394 -5877 2399 -5873
rect 2396 -5884 2399 -5877
rect 2452 -5884 2455 -5867
rect 2513 -5874 2516 -5863
rect 2594 -5866 2600 -5862
rect 2511 -5878 2516 -5874
rect 2513 -5884 2516 -5878
rect 2597 -5884 2600 -5866
rect 2620 -5868 2623 -5853
rect 2618 -5872 2623 -5868
rect 2620 -5884 2623 -5872
rect 2643 -5876 2646 -5853
rect 2641 -5880 2646 -5876
rect 2643 -5884 2646 -5880
rect 2666 -5884 2669 -5853
rect 2722 -5863 2725 -5853
rect 2787 -5858 2790 -5855
rect 2720 -5867 2725 -5863
rect 2722 -5884 2725 -5867
rect 2787 -5875 2790 -5864
rect 2877 -5873 2880 -5853
rect 2785 -5879 2790 -5875
rect 2875 -5877 2880 -5873
rect 2787 -5885 2790 -5879
rect 2877 -5884 2880 -5877
rect 2900 -5884 2903 -5853
rect 2923 -5884 2926 -5853
rect 2946 -5884 2949 -5853
rect 2969 -5884 2972 -5853
rect 3025 -5863 3028 -5853
rect 3023 -5867 3028 -5863
rect 3025 -5884 3028 -5867
rect 2102 -5897 2105 -5890
rect 2149 -5893 2152 -5889
rect 2172 -5905 2175 -5889
rect 2228 -5893 2231 -5889
rect 2285 -5896 2288 -5889
rect 2350 -5893 2353 -5889
rect 2373 -5893 2376 -5889
rect 2396 -5893 2399 -5889
rect 2452 -5893 2455 -5889
rect 2513 -5896 2516 -5889
rect 2597 -5893 2600 -5889
rect 2620 -5893 2623 -5889
rect 2643 -5893 2646 -5889
rect 2149 -5908 2175 -5905
rect 2666 -5908 2669 -5889
rect 2722 -5893 2725 -5889
rect 2787 -5897 2790 -5890
rect 2877 -5893 2880 -5889
rect 2067 -5971 2117 -5968
rect 2067 -6066 2070 -5971
rect 2091 -5990 2094 -5986
rect 2114 -5990 2117 -5971
rect 2145 -5990 2148 -5909
rect 2900 -5917 2903 -5889
rect 2923 -5917 2926 -5889
rect 2946 -5918 2949 -5889
rect 2969 -5917 2972 -5889
rect 3025 -5893 3028 -5889
rect 2168 -5990 2171 -5951
rect 2225 -5995 2228 -5992
rect 2091 -6035 2094 -5996
rect 2114 -6002 2117 -5996
rect 2145 -6014 2148 -5996
rect 2168 -6014 2171 -5996
rect 2225 -6012 2228 -6001
rect 2143 -6018 2148 -6014
rect 2161 -6018 2171 -6014
rect 2091 -6038 2117 -6035
rect 2091 -6045 2094 -6041
rect 2114 -6045 2117 -6038
rect 2145 -6045 2148 -6018
rect 2168 -6045 2171 -6018
rect 2223 -6016 2228 -6012
rect 2091 -6066 2094 -6049
rect 2114 -6053 2117 -6049
rect 2145 -6052 2148 -6049
rect 2168 -6051 2171 -6049
rect 2156 -6053 2171 -6051
rect 2114 -6055 2136 -6053
rect 2134 -6057 2136 -6055
rect 2156 -6057 2158 -6053
rect 2134 -6059 2158 -6057
rect 2187 -6066 2190 -6018
rect 2225 -6022 2228 -6016
rect 2225 -6034 2228 -6027
rect 2067 -6069 2190 -6066
rect -1598 -6149 -1548 -6146
rect -1598 -6244 -1595 -6149
rect -1574 -6168 -1571 -6164
rect -1551 -6168 -1548 -6149
rect -1520 -6168 -1517 -6081
rect 2157 -6083 2160 -6080
rect 2003 -6086 2160 -6083
rect 2003 -6087 2147 -6086
rect -1497 -6168 -1494 -6111
rect -808 -6149 -758 -6146
rect -1574 -6213 -1571 -6174
rect -1551 -6180 -1548 -6174
rect -1520 -6192 -1517 -6174
rect -1522 -6196 -1517 -6192
rect -1574 -6216 -1548 -6213
rect -1574 -6223 -1571 -6219
rect -1551 -6223 -1548 -6216
rect -1520 -6223 -1517 -6196
rect -1497 -6223 -1494 -6174
rect -1574 -6244 -1571 -6227
rect -1551 -6231 -1548 -6227
rect -1520 -6230 -1517 -6227
rect -1497 -6229 -1494 -6227
rect -1509 -6231 -1494 -6229
rect -1551 -6233 -1529 -6231
rect -1531 -6235 -1529 -6233
rect -1509 -6235 -1507 -6231
rect -1531 -6237 -1507 -6235
rect -1478 -6244 -1475 -6196
rect -1598 -6247 -1475 -6244
rect -808 -6244 -805 -6149
rect -784 -6168 -781 -6164
rect -761 -6168 -758 -6149
rect -730 -6168 -727 -6094
rect -707 -6168 -704 -6111
rect 174 -6149 224 -6146
rect -784 -6213 -781 -6174
rect -761 -6180 -758 -6174
rect -730 -6192 -727 -6174
rect -732 -6196 -727 -6192
rect -784 -6216 -758 -6213
rect -784 -6223 -781 -6219
rect -761 -6223 -758 -6216
rect -730 -6223 -727 -6196
rect -707 -6223 -704 -6174
rect -784 -6244 -781 -6227
rect -761 -6231 -758 -6227
rect -730 -6230 -727 -6227
rect -707 -6229 -704 -6227
rect -719 -6231 -704 -6229
rect -761 -6233 -739 -6231
rect -741 -6235 -739 -6233
rect -719 -6235 -717 -6231
rect -741 -6237 -717 -6235
rect -688 -6244 -685 -6196
rect -808 -6247 -685 -6244
rect 174 -6244 177 -6149
rect 198 -6168 201 -6164
rect 221 -6168 224 -6149
rect 252 -6168 255 -6099
rect 275 -6168 278 -6111
rect 1058 -6149 1108 -6146
rect 198 -6213 201 -6174
rect 221 -6180 224 -6174
rect 252 -6192 255 -6174
rect 250 -6196 255 -6192
rect 198 -6216 224 -6213
rect 198 -6223 201 -6219
rect 221 -6223 224 -6216
rect 252 -6223 255 -6196
rect 275 -6223 278 -6174
rect 198 -6244 201 -6227
rect 221 -6231 224 -6227
rect 252 -6230 255 -6227
rect 275 -6229 278 -6227
rect 263 -6231 278 -6229
rect 221 -6233 243 -6231
rect 241 -6235 243 -6233
rect 263 -6235 265 -6231
rect 241 -6237 265 -6235
rect 294 -6244 297 -6196
rect 174 -6247 297 -6244
rect 1058 -6244 1061 -6149
rect 1082 -6168 1085 -6164
rect 1105 -6168 1108 -6149
rect 1136 -6168 1139 -6101
rect 1159 -6168 1162 -6111
rect 2066 -6116 2116 -6113
rect 1082 -6213 1085 -6174
rect 1105 -6180 1108 -6174
rect 1136 -6192 1139 -6174
rect 1134 -6196 1139 -6192
rect 1082 -6216 1108 -6213
rect 1082 -6223 1085 -6219
rect 1105 -6223 1108 -6216
rect 1136 -6223 1139 -6196
rect 1159 -6223 1162 -6174
rect 1082 -6244 1085 -6227
rect 1105 -6231 1108 -6227
rect 1136 -6230 1139 -6227
rect 1159 -6229 1162 -6227
rect 1147 -6231 1162 -6229
rect 1105 -6233 1127 -6231
rect 1125 -6235 1127 -6233
rect 1147 -6235 1149 -6231
rect 1125 -6237 1149 -6235
rect 1178 -6244 1181 -6196
rect 2066 -6211 2069 -6116
rect 2090 -6135 2093 -6131
rect 2113 -6135 2116 -6116
rect 2144 -6135 2147 -6087
rect 2167 -6135 2170 -6089
rect 2224 -6140 2227 -6137
rect 2090 -6159 2093 -6141
rect 2113 -6147 2116 -6141
rect 2144 -6159 2147 -6141
rect 2167 -6159 2170 -6141
rect 2224 -6157 2227 -6146
rect 2079 -6163 2093 -6159
rect 2142 -6163 2147 -6159
rect 2160 -6163 2170 -6159
rect 2090 -6180 2093 -6163
rect 2090 -6183 2116 -6180
rect 2090 -6190 2093 -6186
rect 2113 -6190 2116 -6183
rect 2144 -6190 2147 -6163
rect 2167 -6190 2170 -6163
rect 2222 -6161 2227 -6157
rect 2090 -6211 2093 -6194
rect 2113 -6198 2116 -6194
rect 2144 -6197 2147 -6194
rect 2167 -6196 2170 -6194
rect 2155 -6198 2170 -6196
rect 2113 -6200 2135 -6198
rect 2133 -6202 2135 -6200
rect 2155 -6202 2157 -6198
rect 2133 -6204 2157 -6202
rect 2186 -6211 2189 -6163
rect 2224 -6167 2227 -6161
rect 2224 -6179 2227 -6172
rect 2066 -6214 2189 -6211
rect 2354 -6222 2357 -6219
rect 2377 -6222 2380 -6219
rect 2400 -6222 2403 -6219
rect 2423 -6222 2426 -6219
rect 2479 -6222 2482 -6219
rect 1058 -6247 1181 -6244
rect 1974 -6248 2147 -6245
rect 2144 -6251 2147 -6248
rect 2066 -6278 2116 -6275
rect 2066 -6373 2069 -6278
rect 2090 -6297 2093 -6293
rect 2113 -6297 2116 -6278
rect 2144 -6297 2147 -6256
rect 2167 -6297 2170 -6232
rect 2354 -6248 2357 -6228
rect 2352 -6252 2357 -6248
rect 2354 -6259 2357 -6252
rect 2377 -6259 2380 -6228
rect 2400 -6259 2403 -6228
rect 2423 -6259 2426 -6228
rect 2479 -6238 2482 -6228
rect 2477 -6242 2482 -6238
rect 2479 -6259 2482 -6242
rect 2354 -6268 2357 -6264
rect 2377 -6279 2380 -6264
rect 2400 -6279 2403 -6264
rect 2423 -6280 2426 -6264
rect 2479 -6268 2482 -6264
rect 2224 -6302 2227 -6299
rect 2090 -6320 2093 -6303
rect 2113 -6309 2116 -6303
rect 2079 -6324 2093 -6320
rect 2144 -6321 2147 -6303
rect 2167 -6321 2170 -6303
rect 2224 -6319 2227 -6308
rect 2090 -6342 2093 -6324
rect 2142 -6325 2147 -6321
rect 2160 -6325 2170 -6321
rect 2090 -6345 2116 -6342
rect 2090 -6352 2093 -6348
rect 2113 -6352 2116 -6345
rect 2144 -6352 2147 -6325
rect 2167 -6352 2170 -6325
rect 2222 -6323 2227 -6319
rect 2090 -6373 2093 -6356
rect 2113 -6360 2116 -6356
rect 2144 -6359 2147 -6356
rect 2167 -6358 2170 -6356
rect 2155 -6360 2170 -6358
rect 2113 -6362 2135 -6360
rect 2133 -6364 2135 -6362
rect 2155 -6364 2157 -6360
rect 2133 -6366 2157 -6364
rect 2186 -6373 2189 -6325
rect 2224 -6329 2227 -6323
rect 2224 -6341 2227 -6334
rect 2066 -6376 2189 -6373
rect -1585 -6460 -1535 -6457
rect -1585 -6555 -1582 -6460
rect -1561 -6479 -1558 -6475
rect -1538 -6479 -1535 -6460
rect -1507 -6479 -1504 -6405
rect -1484 -6479 -1481 -6416
rect -1430 -6459 -1380 -6456
rect -1561 -6524 -1558 -6485
rect -1538 -6491 -1535 -6485
rect -1507 -6503 -1504 -6485
rect -1509 -6507 -1504 -6503
rect -1561 -6527 -1535 -6524
rect -1561 -6534 -1558 -6530
rect -1538 -6534 -1535 -6527
rect -1507 -6534 -1504 -6507
rect -1484 -6534 -1481 -6485
rect -1561 -6555 -1558 -6538
rect -1538 -6542 -1535 -6538
rect -1507 -6541 -1504 -6538
rect -1484 -6540 -1481 -6538
rect -1496 -6541 -1481 -6540
rect -1496 -6542 -1485 -6541
rect -1538 -6544 -1516 -6542
rect -1518 -6546 -1516 -6544
rect -1496 -6546 -1494 -6542
rect -1518 -6548 -1494 -6546
rect -1465 -6555 -1460 -6507
rect -1585 -6558 -1460 -6555
rect -1430 -6554 -1427 -6459
rect -1406 -6478 -1403 -6474
rect -1383 -6478 -1380 -6459
rect -1352 -6478 -1349 -6474
rect -1329 -6478 -1326 -6450
rect -784 -6458 -734 -6455
rect -1406 -6523 -1403 -6484
rect -1383 -6490 -1380 -6484
rect -1352 -6502 -1349 -6484
rect -1354 -6506 -1349 -6502
rect -1406 -6526 -1380 -6523
rect -1406 -6533 -1403 -6529
rect -1383 -6533 -1380 -6526
rect -1352 -6533 -1349 -6506
rect -1329 -6533 -1326 -6484
rect -1406 -6554 -1403 -6537
rect -1383 -6541 -1380 -6537
rect -1352 -6540 -1349 -6537
rect -1329 -6539 -1326 -6537
rect -1341 -6540 -1326 -6539
rect -1341 -6541 -1330 -6540
rect -1383 -6543 -1361 -6541
rect -1363 -6545 -1361 -6543
rect -1341 -6545 -1339 -6541
rect -1363 -6547 -1339 -6545
rect -1310 -6554 -1305 -6506
rect -1430 -6557 -1305 -6554
rect -784 -6553 -781 -6458
rect -760 -6477 -757 -6473
rect -737 -6477 -734 -6458
rect -706 -6477 -703 -6394
rect 1946 -6400 2145 -6397
rect -683 -6477 -680 -6407
rect -629 -6457 -579 -6454
rect -760 -6522 -757 -6483
rect -737 -6489 -734 -6483
rect -706 -6501 -703 -6483
rect -708 -6505 -703 -6501
rect -760 -6525 -734 -6522
rect -760 -6532 -757 -6528
rect -737 -6532 -734 -6525
rect -706 -6532 -703 -6505
rect -683 -6532 -680 -6483
rect -760 -6553 -757 -6536
rect -737 -6540 -734 -6536
rect -706 -6539 -703 -6536
rect -683 -6538 -680 -6536
rect -695 -6539 -680 -6538
rect -695 -6540 -684 -6539
rect -737 -6542 -715 -6540
rect -717 -6544 -715 -6542
rect -695 -6544 -693 -6540
rect -717 -6546 -693 -6544
rect -664 -6553 -659 -6505
rect -784 -6556 -659 -6553
rect -629 -6552 -626 -6457
rect -605 -6476 -602 -6472
rect -582 -6476 -579 -6457
rect -551 -6476 -548 -6472
rect -528 -6476 -525 -6454
rect 119 -6458 169 -6455
rect -605 -6521 -602 -6482
rect -582 -6488 -579 -6482
rect -551 -6500 -548 -6482
rect -553 -6504 -548 -6500
rect -605 -6524 -579 -6521
rect -605 -6531 -602 -6527
rect -582 -6531 -579 -6524
rect -551 -6531 -548 -6504
rect -528 -6531 -525 -6482
rect -605 -6552 -602 -6535
rect -582 -6539 -579 -6535
rect -551 -6538 -548 -6535
rect -528 -6537 -525 -6535
rect -540 -6538 -525 -6537
rect -540 -6539 -529 -6538
rect -582 -6541 -560 -6539
rect -562 -6543 -560 -6541
rect -540 -6543 -538 -6539
rect -562 -6545 -538 -6543
rect -509 -6552 -504 -6504
rect -629 -6555 -504 -6552
rect 119 -6553 122 -6458
rect 143 -6477 146 -6473
rect 166 -6477 169 -6458
rect 197 -6477 200 -6404
rect 220 -6477 223 -6407
rect 274 -6457 324 -6454
rect 143 -6522 146 -6483
rect 166 -6489 169 -6483
rect 197 -6501 200 -6483
rect 195 -6505 200 -6501
rect 143 -6525 169 -6522
rect 143 -6532 146 -6528
rect 166 -6532 169 -6525
rect 197 -6532 200 -6505
rect 220 -6532 223 -6483
rect 143 -6553 146 -6536
rect 166 -6540 169 -6536
rect 197 -6539 200 -6536
rect 220 -6538 223 -6536
rect 208 -6539 223 -6538
rect 208 -6540 219 -6539
rect 166 -6542 188 -6540
rect 186 -6544 188 -6542
rect 208 -6544 210 -6540
rect 186 -6546 210 -6544
rect 239 -6553 244 -6505
rect 119 -6556 244 -6553
rect 274 -6552 277 -6457
rect 298 -6476 301 -6472
rect 321 -6476 324 -6457
rect 352 -6476 355 -6472
rect 375 -6476 378 -6456
rect 987 -6457 1037 -6454
rect 298 -6521 301 -6482
rect 321 -6488 324 -6482
rect 352 -6500 355 -6482
rect 350 -6504 355 -6500
rect 298 -6524 324 -6521
rect 298 -6531 301 -6527
rect 321 -6531 324 -6524
rect 352 -6531 355 -6504
rect 375 -6531 378 -6482
rect 298 -6552 301 -6535
rect 321 -6539 324 -6535
rect 352 -6538 355 -6535
rect 375 -6537 378 -6535
rect 363 -6538 378 -6537
rect 363 -6539 374 -6538
rect 321 -6541 343 -6539
rect 341 -6543 343 -6541
rect 363 -6543 365 -6539
rect 341 -6545 365 -6543
rect 394 -6552 399 -6504
rect 274 -6555 399 -6552
rect 987 -6552 990 -6457
rect 1011 -6476 1014 -6472
rect 1034 -6476 1037 -6457
rect 1065 -6476 1068 -6400
rect 1088 -6476 1091 -6407
rect 2067 -6432 2117 -6429
rect 1142 -6456 1192 -6453
rect 1011 -6521 1014 -6482
rect 1034 -6488 1037 -6482
rect 1065 -6500 1068 -6482
rect 1063 -6504 1068 -6500
rect 1011 -6524 1037 -6521
rect 1011 -6531 1014 -6527
rect 1034 -6531 1037 -6524
rect 1065 -6531 1068 -6504
rect 1088 -6531 1091 -6482
rect 1011 -6552 1014 -6535
rect 1034 -6539 1037 -6535
rect 1065 -6538 1068 -6535
rect 1088 -6537 1091 -6535
rect 1076 -6538 1091 -6537
rect 1076 -6539 1087 -6538
rect 1034 -6541 1056 -6539
rect 1054 -6543 1056 -6541
rect 1076 -6543 1078 -6539
rect 1054 -6545 1078 -6543
rect 1107 -6552 1112 -6504
rect 987 -6555 1112 -6552
rect 1142 -6551 1145 -6456
rect 1166 -6475 1169 -6471
rect 1189 -6475 1192 -6456
rect 1220 -6475 1223 -6471
rect 1243 -6475 1246 -6456
rect 1166 -6520 1169 -6481
rect 1189 -6487 1192 -6481
rect 1220 -6499 1223 -6481
rect 1218 -6503 1223 -6499
rect 1166 -6523 1192 -6520
rect 1166 -6530 1169 -6526
rect 1189 -6530 1192 -6523
rect 1220 -6530 1223 -6503
rect 1243 -6530 1246 -6481
rect 1166 -6551 1169 -6534
rect 1189 -6538 1192 -6534
rect 1220 -6537 1223 -6534
rect 1243 -6536 1246 -6534
rect 1231 -6537 1246 -6536
rect 1231 -6538 1242 -6537
rect 1189 -6540 1211 -6538
rect 1209 -6542 1211 -6540
rect 1231 -6542 1233 -6538
rect 1209 -6544 1233 -6542
rect 1262 -6551 1267 -6503
rect 2067 -6527 2070 -6432
rect 2091 -6451 2094 -6447
rect 2114 -6451 2117 -6432
rect 2145 -6451 2148 -6400
rect 2168 -6451 2171 -6410
rect 2225 -6456 2228 -6453
rect 2091 -6474 2094 -6457
rect 2114 -6463 2117 -6457
rect 2080 -6478 2094 -6474
rect 2145 -6475 2148 -6457
rect 2168 -6475 2171 -6457
rect 2225 -6473 2228 -6462
rect 2091 -6496 2094 -6478
rect 2143 -6479 2148 -6475
rect 2161 -6479 2171 -6475
rect 2091 -6499 2117 -6496
rect 2091 -6506 2094 -6502
rect 2114 -6506 2117 -6499
rect 2145 -6506 2148 -6479
rect 2168 -6506 2171 -6479
rect 2223 -6477 2228 -6473
rect 2091 -6527 2094 -6510
rect 2114 -6514 2117 -6510
rect 2145 -6513 2148 -6510
rect 2168 -6512 2171 -6510
rect 2156 -6514 2171 -6512
rect 2114 -6516 2136 -6514
rect 2134 -6518 2136 -6516
rect 2156 -6518 2158 -6514
rect 2134 -6520 2158 -6518
rect 2187 -6527 2190 -6479
rect 2225 -6483 2228 -6477
rect 2225 -6495 2228 -6488
rect 2067 -6530 2190 -6527
rect 1142 -6554 1267 -6551
rect -1667 -6630 -1664 -6627
rect -1644 -6630 -1641 -6627
rect -1606 -6630 -1603 -6627
rect -1527 -6629 -1524 -6626
rect -1504 -6629 -1501 -6626
rect -1466 -6629 -1463 -6626
rect -1382 -6628 -1379 -6625
rect -1359 -6628 -1356 -6625
rect -1321 -6628 -1318 -6625
rect -1221 -6631 -1218 -6627
rect -1198 -6631 -1195 -6627
rect -1175 -6631 -1172 -6627
rect -1152 -6631 -1149 -6627
rect -866 -6628 -863 -6625
rect -843 -6628 -840 -6625
rect -805 -6628 -802 -6625
rect -726 -6627 -723 -6624
rect -703 -6627 -700 -6624
rect -665 -6627 -662 -6624
rect -581 -6626 -578 -6623
rect -558 -6626 -555 -6623
rect -520 -6626 -517 -6623
rect -1667 -6647 -1664 -6636
rect -1669 -6651 -1664 -6647
rect -1667 -6667 -1664 -6651
rect -1644 -6656 -1641 -6636
rect -1606 -6646 -1603 -6636
rect -1527 -6646 -1524 -6635
rect -1608 -6650 -1603 -6646
rect -1529 -6650 -1524 -6646
rect -1646 -6660 -1641 -6656
rect -1644 -6667 -1641 -6660
rect -1606 -6667 -1603 -6650
rect -1527 -6666 -1524 -6650
rect -1504 -6655 -1501 -6635
rect -1466 -6645 -1463 -6635
rect -1382 -6645 -1379 -6634
rect -1468 -6649 -1463 -6645
rect -1384 -6649 -1379 -6645
rect -1506 -6659 -1501 -6655
rect -1504 -6666 -1501 -6659
rect -1466 -6666 -1463 -6649
rect -1382 -6665 -1379 -6649
rect -1359 -6654 -1356 -6634
rect -1321 -6644 -1318 -6634
rect -420 -6629 -417 -6625
rect -397 -6629 -394 -6625
rect -374 -6629 -371 -6625
rect -351 -6629 -348 -6625
rect 37 -6628 40 -6625
rect 60 -6628 63 -6625
rect 98 -6628 101 -6625
rect 177 -6627 180 -6624
rect 200 -6627 203 -6624
rect 238 -6627 241 -6624
rect 322 -6626 325 -6623
rect 345 -6626 348 -6623
rect 383 -6626 386 -6623
rect -1323 -6648 -1318 -6644
rect -1361 -6658 -1356 -6654
rect -1359 -6665 -1356 -6658
rect -1321 -6665 -1318 -6648
rect -1221 -6660 -1218 -6637
rect -1198 -6660 -1195 -6637
rect -1175 -6660 -1172 -6637
rect -1152 -6649 -1149 -6637
rect -866 -6645 -863 -6634
rect -868 -6649 -863 -6645
rect -1154 -6653 -1149 -6649
rect -1152 -6660 -1149 -6653
rect -866 -6665 -863 -6649
rect -843 -6654 -840 -6634
rect -805 -6644 -802 -6634
rect -726 -6644 -723 -6633
rect -807 -6648 -802 -6644
rect -728 -6648 -723 -6644
rect -845 -6658 -840 -6654
rect -843 -6665 -840 -6658
rect -805 -6665 -802 -6648
rect -726 -6664 -723 -6648
rect -703 -6653 -700 -6633
rect -665 -6643 -662 -6633
rect -581 -6643 -578 -6632
rect -667 -6647 -662 -6643
rect -583 -6647 -578 -6643
rect -705 -6657 -700 -6653
rect -703 -6664 -700 -6657
rect -665 -6664 -662 -6647
rect -581 -6663 -578 -6647
rect -558 -6652 -555 -6632
rect -520 -6642 -517 -6632
rect 483 -6629 486 -6625
rect 506 -6629 509 -6625
rect 529 -6629 532 -6625
rect 552 -6629 555 -6625
rect 905 -6627 908 -6624
rect 928 -6627 931 -6624
rect 966 -6627 969 -6624
rect 1045 -6626 1048 -6623
rect 1068 -6626 1071 -6623
rect 1106 -6626 1109 -6623
rect 1190 -6625 1193 -6622
rect 1213 -6625 1216 -6622
rect 1251 -6625 1254 -6622
rect -522 -6646 -517 -6642
rect -560 -6656 -555 -6652
rect -558 -6663 -555 -6656
rect -520 -6663 -517 -6646
rect -420 -6658 -417 -6635
rect -397 -6658 -394 -6635
rect -374 -6658 -371 -6635
rect -351 -6647 -348 -6635
rect 37 -6645 40 -6634
rect -353 -6651 -348 -6647
rect 35 -6649 40 -6645
rect -351 -6658 -348 -6651
rect -1221 -6669 -1218 -6665
rect -1667 -6676 -1664 -6672
rect -1644 -6676 -1641 -6672
rect -1606 -6676 -1603 -6672
rect -1527 -6675 -1524 -6671
rect -1504 -6675 -1501 -6671
rect -1466 -6675 -1463 -6671
rect -1382 -6674 -1379 -6670
rect -1359 -6674 -1356 -6670
rect -1321 -6674 -1318 -6670
rect -1198 -6681 -1195 -6665
rect -1175 -6690 -1172 -6665
rect -1152 -6669 -1149 -6665
rect -420 -6667 -417 -6663
rect -866 -6674 -863 -6670
rect -843 -6674 -840 -6670
rect -805 -6674 -802 -6670
rect -726 -6673 -723 -6669
rect -703 -6673 -700 -6669
rect -665 -6673 -662 -6669
rect -581 -6672 -578 -6668
rect -558 -6672 -555 -6668
rect -520 -6672 -517 -6668
rect -397 -6679 -394 -6663
rect -374 -6688 -371 -6663
rect -351 -6667 -348 -6663
rect 37 -6665 40 -6649
rect 60 -6654 63 -6634
rect 98 -6644 101 -6634
rect 177 -6644 180 -6633
rect 96 -6648 101 -6644
rect 175 -6648 180 -6644
rect 58 -6658 63 -6654
rect 60 -6665 63 -6658
rect 98 -6665 101 -6648
rect 177 -6664 180 -6648
rect 200 -6653 203 -6633
rect 238 -6643 241 -6633
rect 322 -6643 325 -6632
rect 236 -6647 241 -6643
rect 320 -6647 325 -6643
rect 198 -6657 203 -6653
rect 200 -6664 203 -6657
rect 238 -6664 241 -6647
rect 322 -6663 325 -6647
rect 345 -6652 348 -6632
rect 383 -6642 386 -6632
rect 1351 -6628 1354 -6624
rect 1374 -6628 1377 -6624
rect 1397 -6628 1400 -6624
rect 1420 -6628 1423 -6624
rect 381 -6646 386 -6642
rect 343 -6656 348 -6652
rect 345 -6663 348 -6656
rect 383 -6663 386 -6646
rect 483 -6658 486 -6635
rect 506 -6658 509 -6635
rect 529 -6658 532 -6635
rect 552 -6647 555 -6635
rect 905 -6644 908 -6633
rect 550 -6651 555 -6647
rect 903 -6648 908 -6644
rect 552 -6658 555 -6651
rect 483 -6667 486 -6663
rect 37 -6674 40 -6670
rect 60 -6674 63 -6670
rect 98 -6674 101 -6670
rect 177 -6673 180 -6669
rect 200 -6673 203 -6669
rect 238 -6673 241 -6669
rect 322 -6672 325 -6668
rect 345 -6672 348 -6668
rect 383 -6672 386 -6668
rect 506 -6679 509 -6663
rect 529 -6688 532 -6663
rect 552 -6667 555 -6663
rect 905 -6664 908 -6648
rect 928 -6653 931 -6633
rect 966 -6643 969 -6633
rect 1045 -6643 1048 -6632
rect 964 -6647 969 -6643
rect 1043 -6647 1048 -6643
rect 926 -6657 931 -6653
rect 928 -6664 931 -6657
rect 966 -6664 969 -6647
rect 1045 -6663 1048 -6647
rect 1068 -6652 1071 -6632
rect 1106 -6642 1109 -6632
rect 1190 -6642 1193 -6631
rect 1104 -6646 1109 -6642
rect 1188 -6646 1193 -6642
rect 1066 -6656 1071 -6652
rect 1068 -6663 1071 -6656
rect 1106 -6663 1109 -6646
rect 1190 -6662 1193 -6646
rect 1213 -6651 1216 -6631
rect 1251 -6641 1254 -6631
rect 1249 -6645 1254 -6641
rect 1211 -6655 1216 -6651
rect 1213 -6662 1216 -6655
rect 1251 -6662 1254 -6645
rect 1351 -6657 1354 -6634
rect 1374 -6657 1377 -6634
rect 1397 -6657 1400 -6634
rect 1420 -6646 1423 -6634
rect 1418 -6650 1423 -6646
rect 1420 -6657 1423 -6650
rect 2143 -6655 2146 -6652
rect 2166 -6655 2169 -6652
rect 2222 -6655 2225 -6652
rect 2352 -6655 2355 -6652
rect 2375 -6655 2378 -6652
rect 2398 -6655 2401 -6574
rect 2644 -6593 2647 -6574
rect 2644 -6597 2697 -6593
rect 2454 -6655 2457 -6652
rect 2598 -6655 2601 -6652
rect 2621 -6655 2624 -6652
rect 2644 -6655 2647 -6597
rect 2667 -6655 2670 -6628
rect 2723 -6655 2726 -6652
rect 2875 -6654 2878 -6651
rect 2898 -6654 2901 -6619
rect 2921 -6654 2924 -6641
rect 2944 -6654 2947 -6640
rect 2967 -6654 2970 -6639
rect 3107 -6648 3110 -6644
rect 3130 -6648 3133 -6644
rect 3153 -6648 3156 -6644
rect 3176 -6648 3179 -6644
rect 3199 -6648 3202 -6644
rect 3023 -6654 3026 -6651
rect 1351 -6666 1354 -6662
rect 905 -6673 908 -6669
rect 928 -6673 931 -6669
rect 966 -6673 969 -6669
rect 1045 -6672 1048 -6668
rect 1068 -6672 1071 -6668
rect 1106 -6672 1109 -6668
rect 1190 -6671 1193 -6667
rect 1213 -6671 1216 -6667
rect 1251 -6671 1254 -6667
rect 1374 -6678 1377 -6662
rect 1397 -6687 1400 -6662
rect 1420 -6666 1423 -6662
rect 2096 -6666 2099 -6663
rect 2096 -6683 2099 -6672
rect 2143 -6681 2146 -6661
rect 2094 -6687 2099 -6683
rect 2141 -6685 2146 -6681
rect 2096 -6693 2099 -6687
rect 2143 -6692 2146 -6685
rect 2166 -6692 2169 -6661
rect 2222 -6671 2225 -6661
rect 2287 -6665 2290 -6662
rect 2352 -6670 2355 -6661
rect 2220 -6675 2225 -6671
rect 2222 -6692 2225 -6675
rect 2287 -6682 2290 -6671
rect 2346 -6674 2355 -6670
rect 2285 -6686 2290 -6682
rect 2287 -6692 2290 -6686
rect 2352 -6692 2355 -6674
rect 2375 -6676 2378 -6661
rect 2373 -6680 2378 -6676
rect 2375 -6692 2378 -6680
rect 2398 -6692 2401 -6661
rect 2454 -6671 2457 -6661
rect 2514 -6665 2517 -6662
rect 2598 -6670 2601 -6661
rect 2452 -6675 2457 -6671
rect 2454 -6692 2457 -6675
rect 2514 -6682 2517 -6671
rect 2595 -6674 2601 -6670
rect 2512 -6686 2517 -6682
rect 2514 -6692 2517 -6686
rect 2598 -6692 2601 -6674
rect 2621 -6692 2624 -6661
rect 2644 -6692 2647 -6661
rect 2667 -6692 2670 -6661
rect 2723 -6671 2726 -6661
rect 2785 -6665 2788 -6662
rect 2721 -6675 2726 -6671
rect 2723 -6692 2726 -6675
rect 2785 -6682 2788 -6671
rect 2875 -6680 2878 -6660
rect 2783 -6686 2788 -6682
rect 2873 -6684 2878 -6680
rect 2785 -6692 2788 -6686
rect 2875 -6691 2878 -6684
rect 2898 -6691 2901 -6660
rect 2921 -6691 2924 -6660
rect 2944 -6691 2947 -6660
rect 2967 -6691 2970 -6660
rect 3023 -6670 3026 -6660
rect 3107 -6668 3110 -6654
rect 3021 -6674 3026 -6670
rect 3099 -6672 3110 -6668
rect 3023 -6691 3026 -6674
rect 3107 -6677 3110 -6672
rect 3130 -6677 3133 -6654
rect 3153 -6677 3156 -6654
rect 3176 -6677 3179 -6654
rect 3199 -6666 3202 -6654
rect 3197 -6670 3202 -6666
rect 3199 -6677 3202 -6670
rect 3107 -6686 3110 -6682
rect 2096 -6705 2099 -6698
rect 2143 -6701 2146 -6697
rect 2166 -6733 2169 -6697
rect 2222 -6701 2225 -6697
rect 2287 -6704 2290 -6697
rect 2352 -6701 2355 -6697
rect 2375 -6701 2378 -6697
rect 2398 -6701 2401 -6697
rect 2454 -6701 2457 -6697
rect 2514 -6704 2517 -6697
rect 2598 -6701 2601 -6697
rect 2621 -6722 2624 -6697
rect 2644 -6701 2647 -6697
rect 2667 -6701 2670 -6697
rect 2723 -6701 2726 -6697
rect 2785 -6704 2788 -6697
rect 2875 -6700 2878 -6696
rect 2898 -6702 2901 -6696
rect 2921 -6702 2924 -6696
rect 2944 -6702 2947 -6696
rect 2967 -6702 2970 -6696
rect 3023 -6700 3026 -6696
rect 3130 -6702 3133 -6682
rect 3153 -6702 3156 -6682
rect 3176 -6698 3179 -6682
rect 3199 -6689 3202 -6682
<< polycontact >>
rect 664 -5032 669 -5028
rect 723 -5030 728 -5026
rect 685 -5041 690 -5037
rect 1114 -5116 1119 -5112
rect 968 -5134 973 -5130
rect 1027 -5132 1032 -5128
rect 989 -5143 994 -5139
rect 1204 -5129 1209 -5125
rect 1265 -5128 1270 -5124
rect 1227 -5138 1232 -5134
rect 1335 -5129 1340 -5125
rect 1396 -5128 1401 -5124
rect 1358 -5138 1363 -5134
rect 1491 -5129 1496 -5125
rect 1552 -5128 1557 -5124
rect 1514 -5138 1519 -5134
rect 1113 -5184 1118 -5180
rect 574 -5301 579 -5297
rect 682 -5301 687 -5297
rect 794 -5301 799 -5297
rect 906 -5301 911 -5297
rect 1017 -5301 1022 -5297
rect 1129 -5301 1134 -5297
rect 1241 -5301 1246 -5297
rect 1353 -5301 1358 -5297
rect 1793 -5299 1798 -5295
rect 1901 -5299 1906 -5295
rect 2013 -5299 2018 -5295
rect 2125 -5299 2130 -5295
rect 2236 -5299 2241 -5295
rect 2348 -5299 2353 -5295
rect 2460 -5299 2465 -5295
rect 2572 -5299 2577 -5295
rect -577 -5308 -572 -5304
rect -469 -5308 -464 -5304
rect -357 -5308 -352 -5304
rect -245 -5308 -240 -5304
rect -134 -5308 -129 -5304
rect -22 -5308 -17 -5304
rect 90 -5308 95 -5304
rect 202 -5308 207 -5304
rect -517 -5347 -512 -5343
rect -409 -5347 -404 -5343
rect -297 -5347 -292 -5343
rect -185 -5347 -180 -5343
rect -74 -5347 -69 -5343
rect 38 -5347 43 -5343
rect 150 -5347 155 -5343
rect 262 -5347 267 -5343
rect 634 -5340 639 -5336
rect 742 -5340 747 -5336
rect 854 -5340 859 -5336
rect 966 -5340 971 -5336
rect 1077 -5340 1082 -5336
rect 1189 -5340 1194 -5336
rect 1301 -5340 1306 -5336
rect 1413 -5340 1418 -5336
rect 1853 -5338 1858 -5334
rect 1961 -5338 1966 -5334
rect 2073 -5338 2078 -5334
rect 2185 -5338 2190 -5334
rect 2296 -5338 2301 -5334
rect 2408 -5338 2413 -5334
rect 2520 -5338 2525 -5334
rect 2632 -5338 2637 -5334
rect 226 -5445 235 -5436
rect 114 -5463 123 -5454
rect 1 -5486 10 -5477
rect -112 -5515 -103 -5506
rect -223 -5536 -214 -5527
rect -335 -5559 -326 -5550
rect -447 -5574 -438 -5565
rect -555 -5586 -546 -5577
rect 1364 -5445 1371 -5438
rect 1248 -5463 1253 -5456
rect 1143 -5487 1151 -5476
rect 1024 -5516 1035 -5506
rect 899 -5537 913 -5525
rect 789 -5558 798 -5549
rect 677 -5574 687 -5567
rect 2595 -5446 2605 -5438
rect 2480 -5463 2490 -5455
rect 2368 -5484 2378 -5476
rect 2258 -5515 2268 -5507
rect 2147 -5534 2157 -5526
rect 2035 -5558 2043 -5551
rect 1923 -5573 1931 -5566
rect 581 -5587 589 -5579
rect 1815 -5585 1823 -5578
rect 2662 -5731 2667 -5727
rect 2576 -5768 2580 -5763
rect 2599 -5768 2603 -5763
rect 2623 -5768 2627 -5763
rect 2646 -5764 2650 -5759
rect -545 -5789 -537 -5781
rect -522 -5789 -514 -5781
rect -405 -5788 -397 -5780
rect -383 -5787 -375 -5779
rect -267 -5788 -259 -5780
rect -244 -5788 -236 -5780
rect -118 -5787 -110 -5779
rect -95 -5787 -87 -5779
rect 2619 -5800 2624 -5793
rect -488 -5831 -483 -5827
rect -349 -5831 -344 -5827
rect -211 -5831 -206 -5827
rect -61 -5831 -56 -5827
rect 2170 -5831 2177 -5825
rect 2371 -5832 2379 -5827
rect 2899 -5831 2904 -5826
rect 2095 -5879 2100 -5875
rect 2142 -5877 2147 -5873
rect 2221 -5867 2226 -5863
rect 2339 -5866 2344 -5862
rect 2278 -5878 2283 -5874
rect 2366 -5872 2371 -5868
rect 2445 -5867 2450 -5863
rect 2389 -5877 2394 -5873
rect 2589 -5866 2594 -5862
rect 2506 -5878 2511 -5874
rect 2613 -5872 2618 -5868
rect 2636 -5880 2641 -5876
rect 2715 -5867 2720 -5863
rect 2780 -5879 2785 -5875
rect 2870 -5877 2875 -5873
rect 3018 -5867 3023 -5863
rect 2144 -5909 2149 -5905
rect 2665 -5912 2670 -5908
rect 2898 -5923 2903 -5917
rect 2922 -5923 2927 -5917
rect 2944 -5924 2949 -5918
rect 2968 -5923 2973 -5917
rect 2167 -5951 2172 -5947
rect 2138 -6018 2143 -6014
rect 2187 -6018 2191 -6013
rect 2218 -6016 2223 -6012
rect -1522 -6081 -1516 -6076
rect 2157 -6080 2162 -6076
rect 1998 -6087 2003 -6083
rect -732 -6094 -726 -6089
rect -1499 -6111 -1492 -6106
rect -1527 -6196 -1522 -6192
rect -1478 -6196 -1474 -6191
rect 251 -6099 256 -6094
rect -710 -6111 -703 -6106
rect -737 -6196 -732 -6192
rect -688 -6196 -684 -6191
rect 1134 -6101 1140 -6096
rect 273 -6111 280 -6106
rect 245 -6196 250 -6192
rect 294 -6196 298 -6191
rect 1159 -6111 1163 -6106
rect 1129 -6196 1134 -6192
rect 1178 -6196 1182 -6191
rect 2167 -6089 2172 -6085
rect 2074 -6163 2079 -6159
rect 2137 -6163 2142 -6159
rect 2186 -6163 2190 -6158
rect 2217 -6161 2222 -6157
rect 2167 -6232 2171 -6227
rect 1970 -6248 1974 -6243
rect 2144 -6256 2148 -6251
rect 2347 -6252 2352 -6248
rect 2472 -6242 2477 -6238
rect 2376 -6283 2381 -6279
rect 2399 -6283 2404 -6279
rect 2422 -6284 2427 -6280
rect 2074 -6324 2079 -6320
rect 2137 -6325 2142 -6321
rect 2186 -6325 2190 -6320
rect 2217 -6323 2222 -6319
rect -708 -6394 -700 -6387
rect -1508 -6405 -1502 -6400
rect -1488 -6416 -1477 -6406
rect -1329 -6450 -1323 -6442
rect -1514 -6507 -1509 -6503
rect -1465 -6507 -1460 -6503
rect -1485 -6545 -1480 -6541
rect -1359 -6506 -1354 -6502
rect -1310 -6506 -1305 -6502
rect -1330 -6544 -1325 -6540
rect -686 -6407 -678 -6400
rect 193 -6404 200 -6397
rect 1064 -6400 1069 -6395
rect 1941 -6400 1946 -6396
rect 2145 -6400 2150 -6396
rect -528 -6454 -523 -6447
rect -713 -6505 -708 -6501
rect -664 -6505 -659 -6501
rect -684 -6543 -679 -6539
rect -558 -6504 -553 -6500
rect -509 -6504 -504 -6500
rect -529 -6542 -524 -6538
rect 218 -6407 227 -6400
rect 190 -6505 195 -6501
rect 239 -6505 244 -6501
rect 219 -6543 224 -6539
rect 375 -6456 380 -6450
rect 345 -6504 350 -6500
rect 394 -6504 399 -6500
rect 374 -6542 379 -6538
rect 1087 -6407 1096 -6400
rect 1058 -6504 1063 -6500
rect 1107 -6504 1112 -6500
rect 1087 -6542 1092 -6538
rect 1243 -6456 1249 -6451
rect 1213 -6503 1218 -6499
rect 1262 -6503 1267 -6499
rect 1242 -6541 1247 -6537
rect 2167 -6410 2172 -6406
rect 2075 -6478 2080 -6474
rect 2138 -6479 2143 -6475
rect 2187 -6479 2191 -6474
rect 2218 -6477 2223 -6473
rect 2397 -6574 2402 -6570
rect 2642 -6574 2647 -6570
rect -1674 -6651 -1669 -6647
rect -1613 -6650 -1608 -6646
rect -1534 -6650 -1529 -6646
rect -1651 -6660 -1646 -6656
rect -1473 -6649 -1468 -6645
rect -1389 -6649 -1384 -6645
rect -1511 -6659 -1506 -6655
rect -1328 -6648 -1323 -6644
rect -1226 -6648 -1221 -6644
rect -1366 -6658 -1361 -6654
rect -873 -6649 -868 -6645
rect -1159 -6653 -1154 -6649
rect -812 -6648 -807 -6644
rect -733 -6648 -728 -6644
rect -850 -6658 -845 -6654
rect -672 -6647 -667 -6643
rect -588 -6647 -583 -6643
rect -710 -6657 -705 -6653
rect -527 -6646 -522 -6642
rect -425 -6646 -420 -6642
rect -565 -6656 -560 -6652
rect -358 -6651 -353 -6647
rect 30 -6649 35 -6645
rect -1198 -6685 -1193 -6681
rect -397 -6683 -392 -6679
rect 91 -6648 96 -6644
rect 170 -6648 175 -6644
rect 53 -6658 58 -6654
rect 231 -6647 236 -6643
rect 315 -6647 320 -6643
rect 193 -6657 198 -6653
rect 376 -6646 381 -6642
rect 478 -6646 483 -6642
rect 338 -6656 343 -6652
rect 545 -6651 550 -6647
rect 898 -6648 903 -6644
rect 506 -6683 511 -6679
rect 959 -6647 964 -6643
rect 1038 -6647 1043 -6643
rect 921 -6657 926 -6653
rect 1099 -6646 1104 -6642
rect 1183 -6646 1188 -6642
rect 1061 -6656 1066 -6652
rect 1244 -6645 1249 -6641
rect 1346 -6645 1351 -6641
rect 1206 -6655 1211 -6651
rect 1413 -6650 1418 -6646
rect 2697 -6597 2702 -6593
rect 2895 -6619 2901 -6615
rect 2664 -6628 2670 -6624
rect 2919 -6641 2925 -6637
rect 2943 -6640 2949 -6636
rect 2965 -6639 2971 -6635
rect 1374 -6682 1379 -6678
rect 2089 -6687 2094 -6683
rect 2136 -6685 2141 -6681
rect -1176 -6694 -1171 -6690
rect -375 -6692 -370 -6688
rect 528 -6692 533 -6688
rect 1396 -6691 1401 -6687
rect 2215 -6675 2220 -6671
rect 2341 -6674 2346 -6670
rect 2280 -6686 2285 -6682
rect 2368 -6680 2373 -6676
rect 2447 -6675 2452 -6671
rect 2590 -6674 2595 -6670
rect 2507 -6686 2512 -6682
rect 2716 -6675 2721 -6671
rect 2778 -6686 2783 -6682
rect 2868 -6684 2873 -6680
rect 3016 -6674 3021 -6670
rect 3093 -6673 3099 -6668
rect 3192 -6670 3197 -6666
rect 3129 -6707 3133 -6702
rect 3153 -6707 3157 -6702
rect 3176 -6703 3180 -6698
rect 2621 -6726 2626 -6722
rect 2165 -6738 2171 -6733
<< metal1 >>
rect 523 -4989 765 -4984
rect 543 -5004 746 -5000
rect -599 -5101 -565 -5100
rect 543 -5101 550 -5004
rect 661 -5010 666 -5004
rect 684 -5010 689 -5004
rect 722 -5010 727 -5004
rect 675 -5026 679 -5016
rect 698 -5026 702 -5016
rect 736 -5026 740 -5016
rect 760 -5026 765 -4989
rect 574 -5032 664 -5028
rect 675 -5030 723 -5026
rect 736 -5030 765 -5026
rect 574 -5075 579 -5032
rect 610 -5041 685 -5037
rect 610 -5062 616 -5041
rect 698 -5047 702 -5030
rect 736 -5047 740 -5030
rect 679 -5052 684 -5047
rect 661 -5061 665 -5052
rect 722 -5060 726 -5052
rect 661 -5064 720 -5061
rect 1096 -5061 1464 -5058
rect 574 -5080 775 -5075
rect 945 -5094 1075 -5091
rect -599 -5107 922 -5101
rect -599 -5108 -565 -5107
rect -599 -5317 -591 -5108
rect 945 -5130 948 -5094
rect 963 -5106 1045 -5102
rect 965 -5112 970 -5106
rect 988 -5112 993 -5106
rect 1026 -5112 1031 -5106
rect 1072 -5112 1075 -5094
rect 1096 -5112 1099 -5061
rect 1153 -5080 1312 -5077
rect 1111 -5089 1137 -5084
rect 1113 -5095 1118 -5089
rect 1127 -5112 1131 -5101
rect 1148 -5112 1151 -5081
rect 1238 -5098 1243 -5090
rect 1196 -5102 1288 -5098
rect 1072 -5116 1114 -5112
rect 1127 -5116 1151 -5112
rect 1203 -5108 1208 -5102
rect 1226 -5108 1231 -5102
rect 1264 -5108 1269 -5102
rect 979 -5128 983 -5118
rect 1002 -5128 1006 -5118
rect 1040 -5128 1044 -5118
rect 1127 -5122 1131 -5116
rect 1148 -5125 1151 -5116
rect 1217 -5124 1221 -5114
rect 1240 -5124 1244 -5114
rect 1278 -5124 1282 -5114
rect 945 -5134 968 -5130
rect 979 -5132 1027 -5128
rect 1040 -5132 1056 -5128
rect 945 -5143 989 -5139
rect 945 -5179 948 -5143
rect 1002 -5149 1006 -5132
rect 1040 -5149 1044 -5132
rect 983 -5154 988 -5149
rect 965 -5162 969 -5154
rect 1026 -5163 1030 -5154
rect 970 -5166 1030 -5163
rect 1053 -5170 1056 -5132
rect 1113 -5135 1117 -5127
rect 1148 -5129 1169 -5125
rect 1174 -5129 1204 -5125
rect 1217 -5128 1265 -5124
rect 1278 -5128 1288 -5124
rect 1308 -5125 1312 -5080
rect 1374 -5098 1379 -5090
rect 1327 -5102 1419 -5098
rect 1334 -5108 1339 -5102
rect 1357 -5108 1362 -5102
rect 1395 -5108 1400 -5102
rect 1348 -5124 1352 -5114
rect 1371 -5124 1375 -5114
rect 1409 -5124 1413 -5114
rect 1105 -5138 1137 -5135
rect 1148 -5138 1227 -5134
rect 1105 -5157 1136 -5152
rect 1112 -5163 1117 -5157
rect 1126 -5180 1130 -5169
rect 1148 -5180 1151 -5138
rect 1240 -5145 1244 -5128
rect 1278 -5145 1282 -5128
rect 1308 -5129 1335 -5125
rect 1348 -5128 1396 -5124
rect 1409 -5128 1419 -5124
rect 1461 -5125 1464 -5061
rect 1512 -5098 1517 -5090
rect 2709 -5098 2717 -5097
rect 1483 -5102 2717 -5098
rect 1490 -5108 1495 -5102
rect 1513 -5108 1518 -5102
rect 1551 -5108 1556 -5102
rect 1504 -5124 1508 -5114
rect 1527 -5124 1531 -5114
rect 1565 -5124 1569 -5114
rect 1332 -5138 1358 -5134
rect 1371 -5145 1375 -5128
rect 1409 -5145 1413 -5128
rect 1461 -5129 1491 -5125
rect 1504 -5128 1552 -5124
rect 1565 -5128 1790 -5124
rect 1221 -5150 1226 -5145
rect 1352 -5150 1357 -5145
rect 1462 -5138 1514 -5134
rect 1203 -5159 1207 -5150
rect 1264 -5159 1268 -5150
rect 1203 -5162 1268 -5159
rect 1334 -5159 1338 -5150
rect 1395 -5159 1399 -5150
rect 1334 -5162 1399 -5159
rect 950 -5184 1113 -5180
rect 1126 -5184 1151 -5180
rect 1231 -5179 1235 -5162
rect 1361 -5179 1365 -5162
rect 1163 -5182 1448 -5179
rect -577 -5196 1052 -5191
rect -577 -5304 -572 -5196
rect 1090 -5211 1093 -5184
rect 1126 -5190 1130 -5184
rect 1148 -5194 1151 -5184
rect 1462 -5194 1465 -5138
rect 1527 -5145 1531 -5128
rect 1565 -5145 1569 -5128
rect 1508 -5150 1513 -5145
rect 1490 -5159 1494 -5150
rect 1551 -5157 1555 -5150
rect 1551 -5159 2674 -5157
rect 1490 -5162 2674 -5159
rect 1526 -5179 1530 -5162
rect 1480 -5182 1530 -5179
rect 1112 -5203 1116 -5195
rect 1148 -5197 1465 -5194
rect 1105 -5206 1135 -5203
rect 1090 -5214 1307 -5211
rect 574 -5225 1169 -5220
rect 574 -5227 580 -5225
rect 574 -5297 579 -5227
rect 1793 -5295 1798 -5174
rect 579 -5301 682 -5298
rect 687 -5301 794 -5298
rect 799 -5301 906 -5298
rect 911 -5301 1017 -5298
rect 1022 -5301 1129 -5298
rect 1134 -5301 1241 -5298
rect 1246 -5301 1353 -5298
rect 1798 -5299 1901 -5296
rect 1906 -5299 2013 -5296
rect 2018 -5299 2125 -5296
rect 2130 -5299 2236 -5296
rect 2241 -5299 2348 -5296
rect 2353 -5299 2460 -5296
rect 2465 -5299 2572 -5296
rect -572 -5308 -469 -5305
rect -464 -5308 -357 -5305
rect -352 -5308 -245 -5305
rect -240 -5308 -134 -5305
rect -129 -5308 -22 -5305
rect -17 -5308 90 -5305
rect 95 -5308 202 -5305
rect 1772 -5309 2655 -5308
rect 1436 -5310 2655 -5309
rect 553 -5312 2655 -5310
rect 553 -5314 1775 -5312
rect 553 -5317 557 -5314
rect -642 -5321 557 -5317
rect 567 -5320 572 -5314
rect 590 -5320 595 -5314
rect 633 -5320 638 -5314
rect 675 -5320 680 -5314
rect 698 -5320 703 -5314
rect 741 -5320 746 -5314
rect 787 -5320 792 -5314
rect 810 -5320 815 -5314
rect 853 -5320 858 -5314
rect 899 -5320 904 -5314
rect 922 -5320 927 -5314
rect 965 -5320 970 -5314
rect 1010 -5320 1015 -5314
rect 1033 -5320 1038 -5314
rect 1076 -5320 1081 -5314
rect 1122 -5320 1127 -5314
rect 1145 -5320 1150 -5314
rect 1188 -5320 1193 -5314
rect 1234 -5320 1239 -5314
rect 1257 -5320 1262 -5314
rect 1300 -5320 1305 -5314
rect 1346 -5320 1351 -5314
rect 1369 -5320 1374 -5314
rect 1412 -5320 1417 -5314
rect 1786 -5318 1791 -5312
rect 1809 -5318 1814 -5312
rect 1852 -5318 1857 -5312
rect 1894 -5318 1899 -5312
rect 1917 -5318 1922 -5312
rect 1960 -5318 1965 -5312
rect 2006 -5318 2011 -5312
rect 2029 -5318 2034 -5312
rect 2072 -5318 2077 -5312
rect 2118 -5318 2123 -5312
rect 2141 -5318 2146 -5312
rect 2184 -5318 2189 -5312
rect 2229 -5318 2234 -5312
rect 2252 -5318 2257 -5312
rect 2295 -5318 2300 -5312
rect 2341 -5318 2346 -5312
rect 2364 -5318 2369 -5312
rect 2407 -5318 2412 -5312
rect 2453 -5318 2458 -5312
rect 2476 -5318 2481 -5312
rect 2519 -5318 2524 -5312
rect 2565 -5318 2570 -5312
rect 2588 -5318 2593 -5312
rect 2631 -5318 2636 -5312
rect -1832 -5795 -1821 -5794
rect -642 -5795 -637 -5321
rect -584 -5327 -579 -5321
rect -561 -5327 -556 -5321
rect -518 -5327 -513 -5321
rect -476 -5327 -471 -5321
rect -453 -5327 -448 -5321
rect -410 -5327 -405 -5321
rect -364 -5327 -359 -5321
rect -341 -5327 -336 -5321
rect -298 -5327 -293 -5321
rect -252 -5327 -247 -5321
rect -229 -5327 -224 -5321
rect -186 -5327 -181 -5321
rect -141 -5327 -136 -5321
rect -118 -5327 -113 -5321
rect -75 -5327 -70 -5321
rect -29 -5327 -24 -5321
rect -6 -5327 -1 -5321
rect 37 -5327 42 -5321
rect 83 -5327 88 -5321
rect 106 -5327 111 -5321
rect 149 -5327 154 -5321
rect 195 -5327 200 -5321
rect 218 -5327 223 -5321
rect 261 -5327 266 -5321
rect -570 -5343 -566 -5333
rect -547 -5343 -543 -5333
rect -504 -5343 -500 -5333
rect -462 -5343 -458 -5333
rect -439 -5343 -435 -5333
rect -396 -5343 -392 -5333
rect -350 -5343 -346 -5333
rect -327 -5343 -323 -5333
rect -284 -5343 -280 -5333
rect -238 -5343 -234 -5333
rect -215 -5343 -211 -5333
rect -172 -5343 -168 -5333
rect -127 -5343 -123 -5333
rect -104 -5343 -100 -5333
rect -61 -5343 -57 -5333
rect -15 -5343 -11 -5333
rect 8 -5343 12 -5333
rect 51 -5343 55 -5333
rect 97 -5343 101 -5333
rect 120 -5343 124 -5333
rect 163 -5343 167 -5333
rect 209 -5343 213 -5333
rect 232 -5343 236 -5333
rect 275 -5343 279 -5333
rect 581 -5336 585 -5326
rect 604 -5336 608 -5326
rect 647 -5336 651 -5326
rect 581 -5340 634 -5336
rect 647 -5340 655 -5336
rect 689 -5336 693 -5326
rect 712 -5336 716 -5326
rect 755 -5336 759 -5326
rect 689 -5340 742 -5336
rect 755 -5340 764 -5336
rect -570 -5347 -517 -5343
rect -504 -5347 -492 -5343
rect -462 -5347 -409 -5343
rect -396 -5347 -383 -5343
rect -350 -5347 -297 -5343
rect -284 -5347 -271 -5343
rect -238 -5347 -185 -5343
rect -172 -5347 -159 -5343
rect -127 -5347 -74 -5343
rect -61 -5347 -48 -5343
rect -15 -5347 38 -5343
rect 51 -5347 64 -5343
rect 97 -5347 150 -5343
rect 163 -5347 176 -5343
rect 209 -5347 262 -5343
rect 275 -5347 288 -5343
rect -547 -5364 -543 -5347
rect -504 -5364 -500 -5347
rect -495 -5362 -492 -5347
rect -566 -5369 -561 -5364
rect -439 -5364 -435 -5347
rect -396 -5364 -392 -5347
rect -386 -5362 -383 -5347
rect -458 -5369 -453 -5364
rect -327 -5364 -323 -5347
rect -284 -5364 -280 -5347
rect -274 -5361 -271 -5347
rect -346 -5369 -341 -5364
rect -215 -5364 -211 -5347
rect -172 -5364 -168 -5347
rect -162 -5361 -159 -5347
rect -234 -5369 -229 -5364
rect -104 -5364 -100 -5347
rect -61 -5364 -57 -5347
rect -51 -5361 -48 -5347
rect -123 -5369 -118 -5364
rect 8 -5364 12 -5347
rect 51 -5364 55 -5347
rect 61 -5362 64 -5347
rect -11 -5369 -6 -5364
rect 120 -5364 124 -5347
rect 163 -5364 167 -5347
rect 173 -5362 176 -5347
rect 101 -5369 106 -5364
rect 232 -5364 236 -5347
rect 275 -5364 279 -5347
rect 285 -5362 288 -5347
rect 604 -5357 608 -5340
rect 647 -5357 651 -5340
rect 712 -5357 716 -5340
rect 755 -5357 759 -5340
rect 801 -5336 805 -5326
rect 824 -5336 828 -5326
rect 867 -5336 871 -5326
rect 801 -5340 854 -5336
rect 867 -5340 875 -5336
rect 824 -5357 828 -5340
rect 867 -5357 871 -5340
rect 913 -5336 917 -5326
rect 936 -5336 940 -5326
rect 979 -5336 983 -5326
rect 1024 -5336 1028 -5326
rect 1047 -5336 1051 -5326
rect 1090 -5336 1094 -5326
rect 913 -5340 966 -5336
rect 979 -5340 986 -5336
rect 936 -5357 940 -5340
rect 979 -5357 983 -5340
rect 1024 -5340 1077 -5336
rect 1090 -5340 1099 -5336
rect 1136 -5336 1140 -5326
rect 1159 -5336 1163 -5326
rect 1202 -5336 1206 -5326
rect 1248 -5336 1252 -5326
rect 1271 -5336 1275 -5326
rect 1314 -5336 1318 -5326
rect 1360 -5336 1364 -5326
rect 1383 -5336 1387 -5326
rect 1426 -5336 1430 -5326
rect 1800 -5334 1804 -5324
rect 1823 -5334 1827 -5324
rect 1866 -5334 1870 -5324
rect 1136 -5340 1189 -5336
rect 1202 -5340 1211 -5336
rect 1047 -5357 1051 -5340
rect 1090 -5357 1094 -5340
rect 1159 -5357 1163 -5340
rect 1202 -5357 1206 -5340
rect 1248 -5340 1301 -5336
rect 1314 -5340 1323 -5336
rect 1271 -5357 1275 -5340
rect 1314 -5357 1318 -5340
rect 1360 -5340 1413 -5336
rect 1426 -5340 1435 -5336
rect 1383 -5357 1387 -5340
rect 1426 -5357 1430 -5340
rect 1800 -5338 1853 -5334
rect 1866 -5338 1875 -5334
rect 1908 -5334 1912 -5324
rect 1931 -5334 1935 -5324
rect 1974 -5334 1978 -5324
rect 2020 -5334 2024 -5324
rect 2043 -5334 2047 -5324
rect 2086 -5334 2090 -5324
rect 2132 -5334 2136 -5324
rect 2155 -5334 2159 -5324
rect 2198 -5334 2202 -5324
rect 2243 -5334 2247 -5324
rect 2266 -5334 2270 -5324
rect 2309 -5334 2313 -5324
rect 2355 -5334 2359 -5324
rect 2378 -5334 2382 -5324
rect 2421 -5334 2425 -5324
rect 2467 -5334 2471 -5324
rect 2490 -5334 2494 -5324
rect 2533 -5334 2537 -5324
rect 2579 -5334 2583 -5324
rect 2602 -5334 2606 -5324
rect 2645 -5334 2649 -5324
rect 1908 -5338 1961 -5334
rect 1974 -5338 1983 -5334
rect 1823 -5355 1827 -5338
rect 1866 -5355 1870 -5338
rect 1931 -5355 1935 -5338
rect 1974 -5355 1978 -5338
rect 2020 -5338 2073 -5334
rect 2086 -5338 2095 -5334
rect 2043 -5355 2047 -5338
rect 2086 -5355 2090 -5338
rect 2132 -5338 2185 -5334
rect 2198 -5338 2208 -5334
rect 2155 -5355 2159 -5338
rect 2198 -5355 2202 -5338
rect 2243 -5338 2296 -5334
rect 2309 -5338 2318 -5334
rect 2266 -5355 2270 -5338
rect 2309 -5355 2313 -5338
rect 2355 -5338 2408 -5334
rect 2421 -5338 2429 -5334
rect 2378 -5355 2382 -5338
rect 2421 -5355 2425 -5338
rect 2467 -5338 2520 -5334
rect 2533 -5338 2542 -5334
rect 2490 -5355 2494 -5338
rect 2533 -5355 2537 -5338
rect 2579 -5338 2632 -5334
rect 2645 -5338 2655 -5334
rect 2602 -5355 2606 -5338
rect 2645 -5355 2649 -5338
rect 585 -5362 590 -5357
rect 693 -5362 698 -5357
rect 805 -5362 810 -5357
rect 917 -5362 922 -5357
rect 1028 -5362 1033 -5357
rect 1140 -5362 1145 -5357
rect 1252 -5362 1257 -5357
rect 1364 -5362 1369 -5357
rect 1804 -5360 1809 -5355
rect 1912 -5360 1917 -5355
rect 2024 -5360 2029 -5355
rect 2136 -5360 2141 -5355
rect 2247 -5360 2252 -5355
rect 2359 -5360 2364 -5355
rect 2471 -5360 2476 -5355
rect 2583 -5360 2588 -5355
rect 213 -5369 218 -5364
rect -584 -5378 -580 -5369
rect -518 -5377 -514 -5369
rect -476 -5377 -472 -5369
rect -518 -5378 -472 -5377
rect -410 -5377 -406 -5369
rect -364 -5377 -360 -5369
rect -410 -5378 -360 -5377
rect -298 -5377 -294 -5369
rect -252 -5377 -248 -5369
rect -298 -5378 -248 -5377
rect -186 -5377 -182 -5369
rect -141 -5377 -137 -5369
rect -186 -5378 -137 -5377
rect -75 -5377 -71 -5369
rect -29 -5377 -25 -5369
rect -75 -5378 -25 -5377
rect 37 -5377 41 -5369
rect 83 -5377 87 -5369
rect 37 -5378 87 -5377
rect 149 -5377 153 -5369
rect 195 -5377 199 -5369
rect 149 -5378 199 -5377
rect 261 -5377 265 -5369
rect 567 -5371 571 -5362
rect 633 -5370 637 -5362
rect 675 -5370 679 -5362
rect 633 -5371 679 -5370
rect 741 -5370 745 -5362
rect 787 -5370 791 -5362
rect 741 -5371 791 -5370
rect 853 -5370 857 -5362
rect 899 -5370 903 -5362
rect 853 -5371 903 -5370
rect 965 -5370 969 -5362
rect 1010 -5370 1014 -5362
rect 965 -5371 1014 -5370
rect 1076 -5370 1080 -5362
rect 1122 -5370 1126 -5362
rect 1076 -5371 1126 -5370
rect 1188 -5370 1192 -5362
rect 1234 -5370 1238 -5362
rect 1188 -5371 1238 -5370
rect 1300 -5370 1304 -5362
rect 1346 -5370 1350 -5362
rect 1300 -5371 1350 -5370
rect 1412 -5370 1416 -5362
rect 1786 -5369 1790 -5360
rect 1852 -5368 1856 -5360
rect 1894 -5368 1898 -5360
rect 1852 -5369 1898 -5368
rect 1960 -5368 1964 -5360
rect 2006 -5368 2010 -5360
rect 1960 -5369 2010 -5368
rect 2072 -5368 2076 -5360
rect 2118 -5368 2122 -5360
rect 2072 -5369 2122 -5368
rect 2184 -5368 2188 -5360
rect 2229 -5368 2233 -5360
rect 2184 -5369 2233 -5368
rect 2295 -5368 2299 -5360
rect 2341 -5368 2345 -5360
rect 2295 -5369 2345 -5368
rect 2407 -5368 2411 -5360
rect 2453 -5368 2457 -5360
rect 2407 -5369 2457 -5368
rect 2519 -5368 2523 -5360
rect 2565 -5368 2569 -5360
rect 2519 -5369 2569 -5368
rect 2631 -5367 2635 -5360
rect 2667 -5367 2673 -5162
rect 2631 -5369 2668 -5367
rect 1730 -5370 2668 -5369
rect 1412 -5371 2668 -5370
rect 567 -5372 2668 -5371
rect 567 -5374 1791 -5372
rect 567 -5377 572 -5374
rect 261 -5378 572 -5377
rect -623 -5381 572 -5378
rect -623 -5780 -618 -5381
rect -510 -5382 -507 -5381
rect 235 -5445 1364 -5439
rect 1371 -5445 2595 -5439
rect 2605 -5445 2612 -5439
rect 123 -5463 1248 -5456
rect 1253 -5463 2480 -5456
rect 796 -5480 1143 -5479
rect 10 -5485 1143 -5480
rect 10 -5486 840 -5485
rect 1823 -5479 2368 -5478
rect 1151 -5484 2368 -5479
rect 1151 -5485 1832 -5484
rect -103 -5514 1024 -5510
rect 841 -5515 1024 -5514
rect 1035 -5511 1915 -5510
rect 2159 -5511 2258 -5510
rect 1035 -5514 2258 -5511
rect 1035 -5515 1824 -5514
rect 1951 -5515 2168 -5514
rect 614 -5529 899 -5528
rect -214 -5535 899 -5529
rect -214 -5536 619 -5535
rect 2021 -5527 2147 -5526
rect 928 -5528 937 -5527
rect 1362 -5528 2147 -5527
rect 913 -5534 2147 -5528
rect 913 -5535 1952 -5534
rect 928 -5536 937 -5535
rect 567 -5553 789 -5552
rect -326 -5558 789 -5553
rect 798 -5558 2035 -5552
rect -326 -5559 624 -5558
rect 566 -5569 625 -5568
rect 566 -5570 677 -5569
rect -438 -5573 677 -5570
rect -438 -5574 625 -5573
rect 1833 -5569 1923 -5568
rect 687 -5572 1923 -5569
rect 687 -5573 1833 -5572
rect -546 -5585 581 -5579
rect 589 -5580 596 -5579
rect 589 -5585 1815 -5580
rect 1823 -5585 1826 -5580
rect 1272 -5602 1344 -5593
rect 1808 -5596 1815 -5595
rect 1312 -5603 1344 -5602
rect -542 -5612 -497 -5608
rect -542 -5781 -539 -5612
rect -403 -5610 -388 -5607
rect -519 -5781 -516 -5637
rect -403 -5780 -400 -5610
rect -269 -5611 -262 -5608
rect -380 -5779 -377 -5661
rect -265 -5780 -262 -5611
rect -157 -5612 -112 -5609
rect -242 -5780 -239 -5686
rect -115 -5779 -112 -5612
rect 526 -5633 1276 -5623
rect 936 -5664 1140 -5655
rect -92 -5779 -89 -5705
rect -1832 -5801 -637 -5795
rect -1832 -5804 -38 -5801
rect -1880 -6271 -1871 -5866
rect -1832 -6110 -1821 -5804
rect -642 -5805 -38 -5804
rect -623 -5859 -618 -5813
rect -550 -5811 -545 -5805
rect -527 -5811 -522 -5805
rect -489 -5811 -484 -5805
rect -411 -5811 -406 -5805
rect -388 -5811 -383 -5805
rect -350 -5811 -345 -5805
rect -273 -5811 -268 -5805
rect -250 -5811 -245 -5805
rect -212 -5811 -207 -5805
rect -123 -5811 -118 -5805
rect -100 -5811 -95 -5805
rect -62 -5811 -57 -5805
rect -536 -5827 -532 -5817
rect -513 -5827 -509 -5817
rect -475 -5827 -471 -5817
rect -397 -5827 -393 -5817
rect -374 -5827 -370 -5817
rect -336 -5827 -332 -5817
rect -259 -5827 -255 -5817
rect -236 -5827 -232 -5817
rect -198 -5827 -194 -5817
rect -109 -5827 -105 -5817
rect -86 -5827 -82 -5817
rect -48 -5827 -44 -5817
rect -536 -5831 -488 -5827
rect -475 -5831 -465 -5827
rect -397 -5831 -349 -5827
rect -336 -5831 -326 -5827
rect -259 -5831 -211 -5827
rect -198 -5831 -188 -5827
rect -109 -5831 -61 -5827
rect -48 -5831 -38 -5827
rect -513 -5848 -509 -5831
rect -475 -5848 -471 -5831
rect -374 -5848 -370 -5831
rect -336 -5848 -332 -5831
rect -236 -5848 -232 -5831
rect -198 -5848 -194 -5831
rect -86 -5848 -82 -5831
rect -48 -5848 -44 -5831
rect -1778 -5862 -618 -5859
rect -532 -5853 -527 -5848
rect -393 -5853 -388 -5848
rect -255 -5853 -250 -5848
rect -105 -5853 -100 -5848
rect -550 -5862 -546 -5853
rect -489 -5862 -485 -5853
rect -411 -5862 -407 -5853
rect -350 -5862 -346 -5853
rect -273 -5862 -269 -5853
rect -212 -5862 -208 -5853
rect -123 -5862 -119 -5853
rect -62 -5862 -58 -5853
rect -1778 -5865 -58 -5862
rect 599 -5880 605 -5679
rect -1522 -5885 605 -5880
rect -1522 -6076 -1516 -5885
rect 704 -5897 712 -5677
rect -732 -5902 712 -5897
rect -732 -6089 -727 -5902
rect 816 -5912 824 -5675
rect 251 -5918 824 -5912
rect 251 -6094 256 -5918
rect 1134 -6096 1140 -5664
rect 1266 -6106 1276 -5633
rect 1328 -5998 1343 -5603
rect 1807 -5601 2094 -5596
rect 1377 -6035 1385 -5605
rect 1754 -5617 1778 -5610
rect 1754 -5626 1760 -5617
rect -1831 -6120 -1822 -6110
rect -1501 -6111 -1499 -6106
rect -1492 -6111 -710 -6106
rect -703 -6111 273 -6106
rect 280 -6111 1159 -6106
rect 1163 -6110 1280 -6106
rect -1831 -6127 1172 -6120
rect -1880 -6679 -1871 -6281
rect -1831 -6440 -1822 -6127
rect -1582 -6143 -1533 -6139
rect -1582 -6168 -1577 -6143
rect -1582 -6223 -1577 -6174
rect -1568 -6158 -1541 -6153
rect -1568 -6168 -1564 -6158
rect -1545 -6168 -1541 -6158
rect -1568 -6223 -1564 -6174
rect -1568 -6262 -1564 -6227
rect -1559 -6223 -1554 -6174
rect -1545 -6223 -1541 -6174
rect -1536 -6192 -1533 -6143
rect -1528 -6151 -1524 -6127
rect -792 -6143 -743 -6139
rect -1528 -6156 -1500 -6151
rect -1528 -6168 -1523 -6156
rect -1505 -6168 -1500 -6156
rect -792 -6168 -787 -6143
rect -1536 -6196 -1527 -6192
rect -1514 -6201 -1510 -6174
rect -1536 -6205 -1510 -6201
rect -1559 -6235 -1554 -6227
rect -1536 -6235 -1533 -6205
rect -1514 -6223 -1510 -6205
rect -1491 -6191 -1487 -6174
rect -1491 -6196 -1478 -6191
rect -1491 -6223 -1487 -6196
rect -1559 -6238 -1533 -6235
rect -792 -6223 -787 -6174
rect -778 -6158 -751 -6153
rect -778 -6168 -774 -6158
rect -755 -6168 -751 -6158
rect -778 -6223 -774 -6174
rect -1528 -6238 -1524 -6227
rect -1505 -6238 -1501 -6227
rect -1528 -6242 -1501 -6238
rect -1528 -6271 -1524 -6242
rect -778 -6262 -774 -6227
rect -769 -6223 -764 -6174
rect -755 -6223 -751 -6174
rect -746 -6192 -743 -6143
rect -738 -6151 -734 -6127
rect 190 -6143 239 -6139
rect -738 -6156 -710 -6151
rect -738 -6168 -733 -6156
rect -715 -6168 -710 -6156
rect 190 -6168 195 -6143
rect -746 -6196 -737 -6192
rect -724 -6201 -720 -6174
rect -746 -6205 -720 -6201
rect -769 -6235 -764 -6227
rect -746 -6235 -743 -6205
rect -724 -6223 -720 -6205
rect -701 -6191 -697 -6174
rect -701 -6196 -688 -6191
rect -701 -6223 -697 -6196
rect -769 -6238 -743 -6235
rect 190 -6223 195 -6174
rect 204 -6158 231 -6153
rect 204 -6168 208 -6158
rect 227 -6168 231 -6158
rect 204 -6223 208 -6174
rect -738 -6238 -734 -6227
rect -715 -6238 -711 -6227
rect -738 -6242 -711 -6238
rect -738 -6270 -734 -6242
rect 204 -6262 208 -6227
rect 213 -6223 218 -6174
rect 227 -6223 231 -6174
rect 236 -6192 239 -6143
rect 244 -6151 248 -6127
rect 1074 -6143 1123 -6139
rect 244 -6156 272 -6151
rect 244 -6168 249 -6156
rect 267 -6168 272 -6156
rect 1074 -6168 1079 -6143
rect 236 -6196 245 -6192
rect 258 -6201 262 -6174
rect 236 -6205 262 -6201
rect 213 -6235 218 -6227
rect 236 -6235 239 -6205
rect 258 -6223 262 -6205
rect 281 -6191 285 -6174
rect 281 -6196 294 -6191
rect 281 -6223 285 -6196
rect 213 -6238 239 -6235
rect 1074 -6223 1079 -6174
rect 1088 -6158 1115 -6153
rect 1088 -6168 1092 -6158
rect 1111 -6168 1115 -6158
rect 1088 -6223 1092 -6174
rect 244 -6238 248 -6227
rect 267 -6238 271 -6227
rect 244 -6242 271 -6238
rect 244 -6270 248 -6242
rect 1088 -6261 1092 -6227
rect 1097 -6223 1102 -6174
rect 1111 -6223 1115 -6174
rect 1120 -6192 1123 -6143
rect 1128 -6151 1132 -6127
rect 1128 -6156 1156 -6151
rect 1128 -6168 1133 -6156
rect 1151 -6168 1156 -6156
rect 1120 -6196 1129 -6192
rect 1142 -6201 1146 -6174
rect 1120 -6205 1146 -6201
rect 1097 -6235 1102 -6227
rect 1120 -6235 1123 -6205
rect 1142 -6223 1146 -6205
rect 1165 -6191 1169 -6174
rect 1165 -6196 1178 -6191
rect 1165 -6223 1169 -6196
rect 1097 -6238 1123 -6235
rect 1128 -6238 1132 -6227
rect 1151 -6238 1155 -6227
rect 1128 -6242 1155 -6238
rect 1128 -6270 1132 -6242
rect -1305 -6271 1179 -6270
rect -1785 -6278 1179 -6271
rect -1569 -6409 -1564 -6295
rect -1508 -6400 -1503 -6308
rect -779 -6401 -774 -6287
rect -708 -6387 -700 -6307
rect 144 -6399 149 -6300
rect -779 -6406 -686 -6401
rect -1569 -6416 -1488 -6409
rect 144 -6404 193 -6399
rect 204 -6401 209 -6286
rect 1020 -6395 1027 -6309
rect 1020 -6400 1064 -6395
rect 1088 -6400 1093 -6290
rect 204 -6407 218 -6401
rect -1353 -6428 1268 -6418
rect -1352 -6440 -1346 -6428
rect -551 -6438 -545 -6428
rect 352 -6438 358 -6428
rect 1220 -6438 1226 -6428
rect -1831 -6445 -1346 -6440
rect -1059 -6442 -1046 -6441
rect -1787 -6608 -1782 -6445
rect -1569 -6454 -1520 -6450
rect -1569 -6479 -1564 -6454
rect -1763 -6575 -1617 -6571
rect -1763 -6679 -1757 -6575
rect -1602 -6588 -1599 -6508
rect -1569 -6534 -1564 -6485
rect -1555 -6469 -1533 -6464
rect -1555 -6479 -1551 -6469
rect -1532 -6479 -1528 -6469
rect -1555 -6534 -1551 -6485
rect -1546 -6534 -1541 -6485
rect -1532 -6534 -1528 -6485
rect -1523 -6503 -1520 -6454
rect -1515 -6462 -1512 -6445
rect -1409 -6453 -1365 -6449
rect -1515 -6467 -1487 -6462
rect -1515 -6479 -1510 -6467
rect -1492 -6479 -1487 -6467
rect -1414 -6478 -1409 -6454
rect -1520 -6507 -1514 -6503
rect -1501 -6512 -1497 -6485
rect -1523 -6516 -1497 -6512
rect -1546 -6546 -1541 -6538
rect -1523 -6546 -1520 -6516
rect -1501 -6534 -1497 -6516
rect -1478 -6503 -1474 -6485
rect -1478 -6507 -1465 -6503
rect -1478 -6534 -1474 -6507
rect -1546 -6549 -1520 -6546
rect -1414 -6533 -1409 -6484
rect -1400 -6468 -1373 -6463
rect -1400 -6478 -1396 -6468
rect -1377 -6478 -1373 -6468
rect -1400 -6533 -1396 -6484
rect -1391 -6533 -1386 -6484
rect -1377 -6533 -1373 -6484
rect -1368 -6502 -1365 -6453
rect -1349 -6461 -1346 -6445
rect -1323 -6450 -1046 -6442
rect -1360 -6466 -1332 -6461
rect -1360 -6478 -1355 -6466
rect -1337 -6478 -1332 -6466
rect -1368 -6506 -1359 -6502
rect -1346 -6511 -1342 -6484
rect -1368 -6515 -1342 -6511
rect -1515 -6549 -1511 -6538
rect -1492 -6549 -1488 -6538
rect -1391 -6545 -1386 -6537
rect -1368 -6545 -1365 -6515
rect -1346 -6533 -1342 -6515
rect -1323 -6502 -1319 -6484
rect -1323 -6506 -1310 -6502
rect -1323 -6533 -1319 -6506
rect -1515 -6553 -1488 -6549
rect -1503 -6571 -1500 -6553
rect -1484 -6559 -1481 -6545
rect -1391 -6548 -1365 -6545
rect -1360 -6548 -1356 -6537
rect -1337 -6548 -1333 -6537
rect -1360 -6552 -1333 -6548
rect -1346 -6571 -1343 -6552
rect -1570 -6575 -1343 -6571
rect -1329 -6580 -1326 -6544
rect -1550 -6584 -1326 -6580
rect -1715 -6592 -1431 -6588
rect -1715 -6647 -1709 -6592
rect -1698 -6599 -1693 -6598
rect -1698 -6602 -1485 -6599
rect -1698 -6603 -1693 -6602
rect -1697 -6635 -1694 -6603
rect -1650 -6620 -1647 -6613
rect -1682 -6624 -1588 -6620
rect -1675 -6630 -1670 -6624
rect -1652 -6630 -1647 -6624
rect -1614 -6630 -1609 -6624
rect -1661 -6646 -1657 -6636
rect -1638 -6646 -1634 -6636
rect -1600 -6646 -1596 -6636
rect -1715 -6651 -1674 -6647
rect -1661 -6650 -1613 -6646
rect -1600 -6650 -1587 -6646
rect -1693 -6660 -1651 -6656
rect -1638 -6667 -1634 -6650
rect -1600 -6667 -1596 -6650
rect -1880 -6681 -1757 -6679
rect -1657 -6672 -1652 -6667
rect -1675 -6681 -1671 -6672
rect -1614 -6681 -1610 -6672
rect -1882 -6684 -1614 -6681
rect -1882 -6690 -1757 -6684
rect -1882 -6803 -1867 -6690
rect -1590 -6702 -1587 -6650
rect -1577 -6655 -1572 -6602
rect -1554 -6646 -1551 -6610
rect -1519 -6619 -1516 -6613
rect -1542 -6623 -1448 -6619
rect -1535 -6629 -1530 -6623
rect -1512 -6629 -1507 -6623
rect -1474 -6629 -1469 -6623
rect -1521 -6645 -1517 -6635
rect -1498 -6645 -1494 -6635
rect -1460 -6645 -1456 -6635
rect -1554 -6650 -1534 -6646
rect -1521 -6649 -1473 -6645
rect -1460 -6649 -1449 -6645
rect -1577 -6659 -1511 -6655
rect -1498 -6666 -1494 -6649
rect -1460 -6666 -1456 -6649
rect -1517 -6671 -1512 -6666
rect -1535 -6680 -1531 -6671
rect -1474 -6679 -1470 -6671
rect -1535 -6681 -1474 -6680
rect -1531 -6683 -1474 -6681
rect -1452 -6690 -1449 -6649
rect -1438 -6654 -1431 -6592
rect -1416 -6645 -1410 -6584
rect -1373 -6612 -1210 -6609
rect -1377 -6618 -1374 -6613
rect -1397 -6622 -1303 -6618
rect -1215 -6619 -1210 -6612
rect -1390 -6628 -1385 -6622
rect -1367 -6628 -1362 -6622
rect -1329 -6628 -1324 -6622
rect -1229 -6623 -1155 -6619
rect -1376 -6644 -1372 -6634
rect -1353 -6644 -1349 -6634
rect -1315 -6644 -1311 -6634
rect -1229 -6631 -1224 -6623
rect -1160 -6631 -1155 -6623
rect -1211 -6637 -1206 -6631
rect -1188 -6637 -1183 -6631
rect -1416 -6649 -1389 -6645
rect -1376 -6648 -1328 -6644
rect -1315 -6648 -1226 -6644
rect -1438 -6658 -1366 -6654
rect -1353 -6665 -1349 -6648
rect -1315 -6665 -1311 -6648
rect -1169 -6649 -1165 -6637
rect -1146 -6649 -1142 -6637
rect -1169 -6653 -1159 -6649
rect -1146 -6653 -1137 -6649
rect -1169 -6654 -1165 -6653
rect -1215 -6657 -1165 -6654
rect -1215 -6660 -1211 -6657
rect -1192 -6660 -1188 -6657
rect -1169 -6660 -1165 -6657
rect -1146 -6660 -1142 -6653
rect -1372 -6670 -1367 -6665
rect -1390 -6678 -1386 -6670
rect -1329 -6678 -1325 -6670
rect -1229 -6672 -1225 -6665
rect -1206 -6672 -1202 -6665
rect -1183 -6672 -1179 -6665
rect -1160 -6672 -1156 -6665
rect -1229 -6673 -1156 -6672
rect -1309 -6676 -1156 -6673
rect -1309 -6678 -1304 -6676
rect -1329 -6679 -1304 -6678
rect -1386 -6682 -1304 -6679
rect -1300 -6685 -1198 -6682
rect -1300 -6690 -1296 -6685
rect -1452 -6694 -1296 -6690
rect -1287 -6694 -1176 -6690
rect -1287 -6702 -1284 -6694
rect -1590 -6707 -1284 -6702
rect -1059 -6746 -1046 -6450
rect -986 -6443 -545 -6438
rect -986 -6606 -981 -6443
rect -768 -6452 -719 -6448
rect -768 -6477 -763 -6452
rect -962 -6573 -816 -6569
rect -962 -6675 -956 -6573
rect -801 -6586 -798 -6506
rect -768 -6532 -763 -6483
rect -754 -6467 -732 -6462
rect -754 -6477 -750 -6467
rect -731 -6477 -727 -6467
rect -754 -6532 -750 -6483
rect -745 -6532 -740 -6483
rect -731 -6532 -727 -6483
rect -722 -6501 -719 -6452
rect -714 -6460 -711 -6443
rect -608 -6451 -564 -6447
rect -714 -6465 -686 -6460
rect -714 -6477 -709 -6465
rect -691 -6477 -686 -6465
rect -613 -6476 -608 -6452
rect -719 -6505 -713 -6501
rect -700 -6510 -696 -6483
rect -722 -6514 -696 -6510
rect -745 -6544 -740 -6536
rect -722 -6544 -719 -6514
rect -700 -6532 -696 -6514
rect -677 -6501 -673 -6483
rect -677 -6505 -664 -6501
rect -677 -6532 -673 -6505
rect -745 -6547 -719 -6544
rect -613 -6531 -608 -6482
rect -599 -6466 -572 -6461
rect -599 -6476 -595 -6466
rect -576 -6476 -572 -6466
rect -599 -6531 -595 -6482
rect -590 -6531 -585 -6482
rect -576 -6531 -572 -6482
rect -567 -6500 -564 -6451
rect -548 -6459 -545 -6443
rect -83 -6443 358 -6438
rect -523 -6454 -217 -6447
rect -559 -6464 -531 -6459
rect -559 -6476 -554 -6464
rect -536 -6476 -531 -6464
rect -567 -6504 -558 -6500
rect -545 -6509 -541 -6482
rect -567 -6513 -541 -6509
rect -714 -6547 -710 -6536
rect -691 -6547 -687 -6536
rect -590 -6543 -585 -6535
rect -567 -6543 -564 -6513
rect -545 -6531 -541 -6513
rect -522 -6500 -518 -6482
rect -522 -6504 -509 -6500
rect -522 -6531 -518 -6504
rect -714 -6551 -687 -6547
rect -702 -6569 -699 -6551
rect -683 -6557 -680 -6543
rect -590 -6546 -564 -6543
rect -559 -6546 -555 -6535
rect -536 -6546 -532 -6535
rect -559 -6550 -532 -6546
rect -545 -6569 -542 -6550
rect -769 -6573 -542 -6569
rect -528 -6578 -525 -6542
rect -749 -6582 -525 -6578
rect -914 -6590 -630 -6586
rect -914 -6645 -908 -6590
rect -897 -6597 -892 -6596
rect -897 -6600 -684 -6597
rect -897 -6601 -892 -6600
rect -896 -6633 -893 -6601
rect -849 -6618 -846 -6611
rect -881 -6622 -787 -6618
rect -874 -6628 -869 -6622
rect -851 -6628 -846 -6622
rect -813 -6628 -808 -6622
rect -860 -6644 -856 -6634
rect -837 -6644 -833 -6634
rect -799 -6644 -795 -6634
rect -914 -6649 -873 -6645
rect -860 -6648 -812 -6644
rect -799 -6648 -786 -6644
rect -892 -6658 -850 -6654
rect -837 -6665 -833 -6648
rect -799 -6665 -795 -6648
rect -856 -6670 -851 -6665
rect -874 -6679 -870 -6670
rect -813 -6679 -809 -6670
rect -953 -6682 -813 -6679
rect -789 -6700 -786 -6648
rect -776 -6653 -771 -6600
rect -753 -6644 -750 -6608
rect -718 -6617 -715 -6611
rect -741 -6621 -647 -6617
rect -734 -6627 -729 -6621
rect -711 -6627 -706 -6621
rect -673 -6627 -668 -6621
rect -720 -6643 -716 -6633
rect -697 -6643 -693 -6633
rect -659 -6643 -655 -6633
rect -753 -6648 -733 -6644
rect -720 -6647 -672 -6643
rect -659 -6647 -648 -6643
rect -776 -6657 -710 -6653
rect -697 -6664 -693 -6647
rect -659 -6664 -655 -6647
rect -716 -6669 -711 -6664
rect -734 -6678 -730 -6669
rect -673 -6677 -669 -6669
rect -734 -6679 -673 -6678
rect -730 -6681 -673 -6679
rect -651 -6688 -648 -6647
rect -637 -6652 -630 -6590
rect -615 -6643 -609 -6582
rect -572 -6610 -409 -6607
rect -576 -6616 -573 -6611
rect -596 -6620 -502 -6616
rect -414 -6617 -409 -6610
rect -589 -6626 -584 -6620
rect -566 -6626 -561 -6620
rect -528 -6626 -523 -6620
rect -428 -6621 -354 -6617
rect -575 -6642 -571 -6632
rect -552 -6642 -548 -6632
rect -514 -6642 -510 -6632
rect -428 -6629 -423 -6621
rect -359 -6629 -354 -6621
rect -410 -6635 -405 -6629
rect -387 -6635 -382 -6629
rect -615 -6647 -588 -6643
rect -575 -6646 -527 -6642
rect -514 -6646 -425 -6642
rect -637 -6656 -565 -6652
rect -552 -6663 -548 -6646
rect -514 -6663 -510 -6646
rect -368 -6647 -364 -6635
rect -345 -6647 -341 -6635
rect -368 -6651 -358 -6647
rect -345 -6651 -330 -6647
rect -368 -6652 -364 -6651
rect -414 -6655 -364 -6652
rect -414 -6658 -410 -6655
rect -391 -6658 -387 -6655
rect -368 -6658 -364 -6655
rect -345 -6658 -341 -6651
rect -571 -6668 -566 -6663
rect -589 -6676 -585 -6668
rect -528 -6676 -524 -6668
rect -428 -6670 -424 -6663
rect -405 -6670 -401 -6663
rect -382 -6670 -378 -6663
rect -359 -6670 -355 -6663
rect -428 -6671 -355 -6670
rect -508 -6674 -355 -6671
rect -508 -6676 -503 -6674
rect -528 -6677 -503 -6676
rect -585 -6680 -503 -6677
rect -499 -6683 -397 -6680
rect -499 -6688 -495 -6683
rect -651 -6692 -495 -6688
rect -486 -6692 -375 -6688
rect -486 -6700 -483 -6692
rect -789 -6705 -483 -6700
rect -337 -6746 -330 -6651
rect -1059 -6759 -330 -6746
rect -231 -6741 -217 -6454
rect -83 -6606 -78 -6443
rect 135 -6452 184 -6448
rect 135 -6477 140 -6452
rect -59 -6573 87 -6569
rect -59 -6678 -53 -6573
rect 102 -6586 105 -6506
rect 135 -6532 140 -6483
rect 149 -6467 171 -6462
rect 149 -6477 153 -6467
rect 172 -6477 176 -6467
rect 149 -6532 153 -6483
rect 158 -6532 163 -6483
rect 172 -6532 176 -6483
rect 181 -6501 184 -6452
rect 189 -6460 192 -6443
rect 295 -6451 339 -6447
rect 189 -6465 217 -6460
rect 189 -6477 194 -6465
rect 212 -6477 217 -6465
rect 290 -6476 295 -6452
rect 184 -6505 190 -6501
rect 203 -6510 207 -6483
rect 181 -6514 207 -6510
rect 158 -6544 163 -6536
rect 181 -6544 184 -6514
rect 203 -6532 207 -6514
rect 226 -6501 230 -6483
rect 226 -6505 239 -6501
rect 226 -6532 230 -6505
rect 158 -6547 184 -6544
rect 290 -6531 295 -6482
rect 304 -6466 331 -6461
rect 304 -6476 308 -6466
rect 327 -6476 331 -6466
rect 304 -6531 308 -6482
rect 313 -6531 318 -6482
rect 327 -6531 331 -6482
rect 336 -6500 339 -6451
rect 355 -6459 358 -6443
rect 785 -6442 1226 -6438
rect 610 -6450 613 -6449
rect 380 -6456 613 -6450
rect 344 -6464 372 -6459
rect 344 -6476 349 -6464
rect 367 -6476 372 -6464
rect 336 -6504 345 -6500
rect 358 -6509 362 -6482
rect 336 -6513 362 -6509
rect 189 -6547 193 -6536
rect 212 -6547 216 -6536
rect 313 -6543 318 -6535
rect 336 -6543 339 -6513
rect 358 -6531 362 -6513
rect 381 -6500 385 -6482
rect 381 -6504 394 -6500
rect 381 -6531 385 -6504
rect 189 -6551 216 -6547
rect 201 -6569 204 -6551
rect 220 -6557 223 -6543
rect 313 -6546 339 -6543
rect 344 -6546 348 -6535
rect 367 -6546 371 -6535
rect 344 -6550 371 -6546
rect 358 -6569 361 -6550
rect 134 -6573 361 -6569
rect 375 -6578 378 -6542
rect 154 -6582 378 -6578
rect -11 -6590 273 -6586
rect -11 -6645 -5 -6590
rect 6 -6597 11 -6596
rect 6 -6600 219 -6597
rect 6 -6601 11 -6600
rect 7 -6633 10 -6601
rect 54 -6618 57 -6611
rect 22 -6622 116 -6618
rect 29 -6628 34 -6622
rect 52 -6628 57 -6622
rect 90 -6628 95 -6622
rect 43 -6644 47 -6634
rect 66 -6644 70 -6634
rect 104 -6644 108 -6634
rect -11 -6649 30 -6645
rect 43 -6648 91 -6644
rect 104 -6648 117 -6644
rect 11 -6658 53 -6654
rect 66 -6665 70 -6648
rect 104 -6665 108 -6648
rect 47 -6670 52 -6665
rect 29 -6679 33 -6670
rect 90 -6679 94 -6670
rect -49 -6682 90 -6679
rect 114 -6700 117 -6648
rect 127 -6653 132 -6600
rect 150 -6644 153 -6608
rect 185 -6617 188 -6611
rect 162 -6621 256 -6617
rect 169 -6627 174 -6621
rect 192 -6627 197 -6621
rect 230 -6627 235 -6621
rect 183 -6643 187 -6633
rect 206 -6643 210 -6633
rect 244 -6643 248 -6633
rect 150 -6648 170 -6644
rect 183 -6647 231 -6643
rect 244 -6647 255 -6643
rect 127 -6657 193 -6653
rect 206 -6664 210 -6647
rect 244 -6664 248 -6647
rect 187 -6669 192 -6664
rect 169 -6678 173 -6669
rect 230 -6677 234 -6669
rect 169 -6679 230 -6678
rect 173 -6681 230 -6679
rect 252 -6688 255 -6647
rect 266 -6652 273 -6590
rect 288 -6643 294 -6582
rect 331 -6610 494 -6607
rect 327 -6616 330 -6611
rect 307 -6620 401 -6616
rect 489 -6617 494 -6610
rect 314 -6626 319 -6620
rect 337 -6626 342 -6620
rect 375 -6626 380 -6620
rect 475 -6621 549 -6617
rect 328 -6642 332 -6632
rect 351 -6642 355 -6632
rect 389 -6642 393 -6632
rect 475 -6629 480 -6621
rect 544 -6629 549 -6621
rect 493 -6635 498 -6629
rect 516 -6635 521 -6629
rect 288 -6647 315 -6643
rect 328 -6646 376 -6642
rect 389 -6646 478 -6642
rect 266 -6656 338 -6652
rect 351 -6663 355 -6646
rect 389 -6663 393 -6646
rect 535 -6647 539 -6635
rect 558 -6647 562 -6635
rect 535 -6651 545 -6647
rect 558 -6651 572 -6647
rect 535 -6652 539 -6651
rect 489 -6655 539 -6652
rect 489 -6658 493 -6655
rect 512 -6658 516 -6655
rect 535 -6658 539 -6655
rect 558 -6658 562 -6651
rect 332 -6668 337 -6663
rect 314 -6676 318 -6668
rect 375 -6676 379 -6668
rect 475 -6670 479 -6663
rect 498 -6670 502 -6663
rect 521 -6670 525 -6663
rect 544 -6670 548 -6663
rect 475 -6671 548 -6670
rect 395 -6674 548 -6671
rect 395 -6676 400 -6674
rect 375 -6677 400 -6676
rect 318 -6680 400 -6677
rect 404 -6683 506 -6680
rect 404 -6688 408 -6683
rect 252 -6692 408 -6688
rect 417 -6692 528 -6688
rect 417 -6700 420 -6692
rect 114 -6705 420 -6700
rect 567 -6741 572 -6651
rect -231 -6756 573 -6741
rect 604 -6746 613 -6456
rect 785 -6605 790 -6442
rect 1003 -6451 1052 -6447
rect 1003 -6476 1008 -6451
rect 809 -6572 955 -6568
rect 809 -6678 815 -6572
rect 970 -6585 973 -6505
rect 1003 -6531 1008 -6482
rect 1017 -6466 1039 -6461
rect 1017 -6476 1021 -6466
rect 1040 -6476 1044 -6466
rect 1017 -6531 1021 -6482
rect 1026 -6531 1031 -6482
rect 1040 -6531 1044 -6482
rect 1049 -6500 1052 -6451
rect 1057 -6459 1060 -6442
rect 1163 -6450 1207 -6446
rect 1057 -6464 1085 -6459
rect 1057 -6476 1062 -6464
rect 1080 -6476 1085 -6464
rect 1158 -6475 1163 -6451
rect 1052 -6504 1058 -6500
rect 1071 -6509 1075 -6482
rect 1049 -6513 1075 -6509
rect 1026 -6543 1031 -6535
rect 1049 -6543 1052 -6513
rect 1071 -6531 1075 -6513
rect 1094 -6500 1098 -6482
rect 1094 -6504 1107 -6500
rect 1094 -6531 1098 -6504
rect 1026 -6546 1052 -6543
rect 1158 -6530 1163 -6481
rect 1172 -6465 1199 -6460
rect 1172 -6475 1176 -6465
rect 1195 -6475 1199 -6465
rect 1172 -6530 1176 -6481
rect 1181 -6530 1186 -6481
rect 1195 -6530 1199 -6481
rect 1204 -6499 1207 -6450
rect 1223 -6458 1226 -6442
rect 1275 -6451 1280 -6110
rect 1249 -6456 1280 -6451
rect 1212 -6463 1240 -6458
rect 1212 -6475 1217 -6463
rect 1235 -6475 1240 -6463
rect 1752 -6473 1760 -5626
rect 1808 -6320 1815 -5601
rect 1843 -5617 2206 -5610
rect 2709 -5697 2717 -5102
rect 2052 -5701 2717 -5697
rect 2732 -5372 2733 -5367
rect 2052 -5702 2574 -5701
rect 1884 -5756 2019 -5750
rect 1984 -6159 1989 -5775
rect 2014 -5931 2019 -5756
rect 2031 -5897 2036 -5754
rect 2052 -5837 2057 -5702
rect 2569 -5709 2574 -5702
rect 2661 -5709 2666 -5701
rect 2732 -5707 2740 -5372
rect 2587 -5715 2592 -5709
rect 2610 -5715 2615 -5709
rect 2633 -5715 2638 -5709
rect 2652 -5727 2656 -5715
rect 2675 -5727 2679 -5715
rect 2695 -5710 2740 -5707
rect 2583 -5731 2662 -5727
rect 2675 -5731 2685 -5727
rect 2583 -5738 2587 -5731
rect 2606 -5738 2610 -5731
rect 2629 -5738 2633 -5731
rect 2652 -5738 2656 -5731
rect 2675 -5738 2679 -5731
rect 2569 -5750 2573 -5743
rect 2592 -5750 2596 -5743
rect 2615 -5750 2619 -5743
rect 2638 -5750 2642 -5743
rect 2661 -5750 2665 -5743
rect 2105 -5751 2665 -5750
rect 2695 -5751 2698 -5710
rect 2105 -5754 2698 -5751
rect 2706 -5755 3049 -5751
rect 2246 -5768 2576 -5763
rect 2172 -5825 2175 -5774
rect 2246 -5825 2250 -5768
rect 2599 -5776 2603 -5768
rect 2706 -5760 2710 -5755
rect 2650 -5764 2710 -5760
rect 2623 -5772 2745 -5768
rect 2470 -5779 2603 -5776
rect 2373 -5827 2376 -5785
rect 2470 -5826 2473 -5779
rect 2548 -5799 2619 -5794
rect 2742 -5829 2745 -5772
rect 2900 -5826 2903 -5772
rect 2052 -5840 3041 -5837
rect 2052 -5841 2468 -5840
rect 2031 -5902 2032 -5897
rect 1984 -6164 1986 -6159
rect 1805 -6325 1954 -6320
rect 1805 -6326 1958 -6325
rect 1751 -6478 1915 -6473
rect 1752 -6480 1760 -6478
rect 1204 -6503 1213 -6499
rect 1226 -6508 1230 -6481
rect 1204 -6512 1230 -6508
rect 1057 -6546 1061 -6535
rect 1080 -6546 1084 -6535
rect 1181 -6542 1186 -6534
rect 1204 -6542 1207 -6512
rect 1226 -6530 1230 -6512
rect 1249 -6499 1253 -6481
rect 1249 -6503 1262 -6499
rect 1249 -6530 1253 -6503
rect 1057 -6550 1084 -6546
rect 1069 -6568 1072 -6550
rect 1088 -6556 1091 -6542
rect 1181 -6545 1207 -6542
rect 1212 -6545 1216 -6534
rect 1235 -6545 1239 -6534
rect 1212 -6549 1239 -6545
rect 1226 -6568 1229 -6549
rect 1002 -6572 1229 -6568
rect 1243 -6577 1246 -6541
rect 1022 -6581 1246 -6577
rect 857 -6589 1141 -6585
rect 857 -6644 863 -6589
rect 874 -6596 879 -6595
rect 874 -6599 1087 -6596
rect 874 -6600 879 -6599
rect 875 -6632 878 -6600
rect 922 -6617 925 -6610
rect 890 -6621 984 -6617
rect 897 -6627 902 -6621
rect 920 -6627 925 -6621
rect 958 -6627 963 -6621
rect 911 -6643 915 -6633
rect 934 -6643 938 -6633
rect 972 -6643 976 -6633
rect 857 -6648 898 -6644
rect 911 -6647 959 -6643
rect 972 -6647 985 -6643
rect 879 -6657 921 -6653
rect 934 -6664 938 -6647
rect 972 -6664 976 -6647
rect 915 -6669 920 -6664
rect 897 -6678 901 -6669
rect 958 -6678 962 -6669
rect 819 -6681 958 -6678
rect 982 -6699 985 -6647
rect 995 -6652 1000 -6599
rect 1018 -6643 1021 -6607
rect 1053 -6616 1056 -6610
rect 1030 -6620 1124 -6616
rect 1037 -6626 1042 -6620
rect 1060 -6626 1065 -6620
rect 1098 -6626 1103 -6620
rect 1051 -6642 1055 -6632
rect 1074 -6642 1078 -6632
rect 1112 -6642 1116 -6632
rect 1018 -6647 1038 -6643
rect 1051 -6646 1099 -6642
rect 1112 -6646 1123 -6642
rect 995 -6656 1061 -6652
rect 1074 -6663 1078 -6646
rect 1112 -6663 1116 -6646
rect 1055 -6668 1060 -6663
rect 1037 -6677 1041 -6668
rect 1098 -6676 1102 -6668
rect 1037 -6678 1098 -6677
rect 1041 -6680 1098 -6678
rect 1120 -6687 1123 -6646
rect 1134 -6651 1141 -6589
rect 1156 -6642 1162 -6581
rect 1199 -6609 1362 -6606
rect 1195 -6615 1198 -6610
rect 1175 -6619 1269 -6615
rect 1357 -6616 1362 -6609
rect 1182 -6625 1187 -6619
rect 1205 -6625 1210 -6619
rect 1243 -6625 1248 -6619
rect 1343 -6620 1417 -6616
rect 1196 -6641 1200 -6631
rect 1219 -6641 1223 -6631
rect 1257 -6641 1261 -6631
rect 1343 -6628 1348 -6620
rect 1412 -6628 1417 -6620
rect 1361 -6634 1366 -6628
rect 1384 -6634 1389 -6628
rect 1156 -6646 1183 -6642
rect 1196 -6645 1244 -6641
rect 1257 -6645 1346 -6641
rect 1134 -6655 1206 -6651
rect 1219 -6662 1223 -6645
rect 1257 -6662 1261 -6645
rect 1403 -6646 1407 -6634
rect 1426 -6646 1430 -6634
rect 1403 -6650 1413 -6646
rect 1426 -6650 1437 -6646
rect 1403 -6651 1407 -6650
rect 1357 -6654 1407 -6651
rect 1357 -6657 1361 -6654
rect 1380 -6657 1384 -6654
rect 1403 -6657 1407 -6654
rect 1426 -6657 1430 -6650
rect 1200 -6667 1205 -6662
rect 1182 -6675 1186 -6667
rect 1243 -6675 1247 -6667
rect 1343 -6669 1347 -6662
rect 1366 -6669 1370 -6662
rect 1389 -6669 1393 -6662
rect 1412 -6669 1416 -6662
rect 1343 -6670 1416 -6669
rect 1263 -6673 1416 -6670
rect 1263 -6675 1268 -6673
rect 1243 -6676 1268 -6675
rect 1186 -6679 1268 -6676
rect 1272 -6682 1374 -6679
rect 1272 -6687 1276 -6682
rect 1120 -6691 1276 -6687
rect 1285 -6691 1396 -6687
rect 1285 -6699 1288 -6691
rect 982 -6704 1288 -6699
rect 1434 -6746 1437 -6650
rect 604 -6756 1438 -6746
rect 604 -6757 793 -6756
rect -1882 -6811 -964 -6803
rect -1874 -6813 -964 -6811
rect -953 -6813 -60 -6803
rect -49 -6813 809 -6803
rect 820 -6813 823 -6803
rect 1941 -6812 1945 -6400
rect 1954 -6804 1958 -6326
rect 1970 -6789 1974 -6248
rect 1986 -6764 1991 -6164
rect 1998 -6748 2003 -6087
rect 2014 -6733 2019 -5936
rect 2022 -6719 2027 -5910
rect 2031 -6076 2036 -5902
rect 2052 -5944 2057 -5841
rect 2087 -5847 2091 -5841
rect 2141 -5847 2146 -5841
rect 2164 -5847 2169 -5841
rect 2220 -5847 2225 -5841
rect 2270 -5846 2275 -5841
rect 2087 -5852 2118 -5847
rect 2094 -5858 2099 -5852
rect 2270 -5851 2301 -5846
rect 2342 -5847 2347 -5841
rect 2365 -5847 2370 -5841
rect 2388 -5847 2393 -5841
rect 2444 -5847 2449 -5841
rect 2498 -5846 2503 -5840
rect 2559 -5841 3041 -5840
rect 2108 -5875 2112 -5864
rect 2155 -5863 2159 -5853
rect 2178 -5863 2182 -5853
rect 2234 -5863 2238 -5853
rect 2277 -5857 2282 -5851
rect 2498 -5851 2529 -5846
rect 2589 -5847 2594 -5841
rect 2612 -5847 2617 -5841
rect 2635 -5847 2640 -5841
rect 2658 -5847 2663 -5841
rect 2714 -5847 2719 -5841
rect 2772 -5847 2776 -5841
rect 2869 -5847 2874 -5841
rect 2892 -5847 2897 -5841
rect 2915 -5847 2920 -5841
rect 2938 -5847 2943 -5841
rect 2961 -5847 2966 -5841
rect 3017 -5847 3022 -5841
rect 2155 -5867 2221 -5863
rect 2234 -5867 2244 -5863
rect 2356 -5862 2360 -5853
rect 2379 -5862 2383 -5853
rect 2402 -5862 2406 -5853
rect 2117 -5875 2142 -5873
rect 2065 -5879 2095 -5875
rect 2108 -5877 2142 -5875
rect 2108 -5879 2121 -5877
rect 2065 -5931 2069 -5879
rect 2108 -5885 2112 -5879
rect 2178 -5884 2182 -5867
rect 2234 -5884 2238 -5867
rect 2291 -5874 2295 -5863
rect 2302 -5866 2339 -5862
rect 2356 -5863 2406 -5862
rect 2458 -5863 2462 -5853
rect 2505 -5857 2510 -5851
rect 2772 -5852 2803 -5847
rect 2356 -5865 2445 -5863
rect 2302 -5874 2305 -5866
rect 2402 -5867 2445 -5865
rect 2458 -5867 2468 -5863
rect 2603 -5862 2607 -5853
rect 2626 -5862 2630 -5853
rect 2649 -5862 2653 -5853
rect 2672 -5862 2676 -5853
rect 2250 -5878 2278 -5874
rect 2291 -5878 2305 -5874
rect 2308 -5872 2366 -5869
rect 2291 -5884 2295 -5878
rect 2308 -5881 2311 -5872
rect 2386 -5875 2389 -5874
rect 2159 -5889 2164 -5884
rect 2300 -5884 2311 -5881
rect 2320 -5878 2389 -5875
rect 2300 -5889 2303 -5884
rect 2094 -5898 2098 -5890
rect 2141 -5898 2145 -5889
rect 2220 -5898 2224 -5889
rect 2277 -5898 2281 -5889
rect 2320 -5890 2323 -5878
rect 2402 -5884 2406 -5867
rect 2458 -5884 2462 -5867
rect 2519 -5874 2523 -5863
rect 2532 -5866 2589 -5862
rect 2603 -5863 2676 -5862
rect 2728 -5863 2732 -5853
rect 2779 -5858 2784 -5852
rect 2603 -5865 2715 -5863
rect 2532 -5874 2536 -5866
rect 2672 -5867 2715 -5865
rect 2728 -5867 2741 -5863
rect 2477 -5878 2506 -5874
rect 2519 -5878 2536 -5874
rect 2539 -5872 2613 -5869
rect 2519 -5884 2523 -5878
rect 2539 -5882 2542 -5872
rect 2314 -5893 2323 -5890
rect 2360 -5889 2365 -5884
rect 2383 -5889 2388 -5884
rect 2528 -5885 2542 -5882
rect 2547 -5880 2636 -5876
rect 2342 -5898 2346 -5889
rect 2444 -5898 2448 -5889
rect 2505 -5898 2509 -5889
rect 2528 -5890 2532 -5885
rect 2547 -5890 2550 -5880
rect 2672 -5884 2676 -5867
rect 2728 -5884 2732 -5867
rect 2793 -5875 2797 -5864
rect 2883 -5863 2887 -5853
rect 2906 -5863 2910 -5853
rect 2929 -5863 2933 -5853
rect 2952 -5863 2956 -5853
rect 2975 -5863 2979 -5853
rect 3031 -5863 3035 -5853
rect 3045 -5863 3049 -5755
rect 2883 -5867 3018 -5863
rect 3031 -5867 3049 -5863
rect 2860 -5875 2870 -5873
rect 2765 -5879 2780 -5875
rect 2793 -5878 2870 -5875
rect 2793 -5879 2861 -5878
rect 2607 -5889 2612 -5884
rect 2630 -5889 2635 -5884
rect 2653 -5889 2658 -5884
rect 2793 -5885 2797 -5879
rect 2975 -5884 2979 -5867
rect 3031 -5884 3035 -5867
rect 2589 -5898 2593 -5889
rect 2714 -5898 2718 -5889
rect 2887 -5889 2892 -5884
rect 2910 -5889 2915 -5884
rect 2933 -5889 2938 -5884
rect 2956 -5889 2961 -5884
rect 2779 -5898 2783 -5890
rect 2869 -5898 2873 -5889
rect 3017 -5898 3021 -5889
rect 2091 -5901 3021 -5898
rect 2718 -5902 2870 -5901
rect 2111 -5908 2144 -5905
rect 2666 -5925 2669 -5912
rect 2065 -5938 2070 -5936
rect 2279 -5932 2471 -5927
rect 2579 -5930 2669 -5925
rect 2065 -5941 2171 -5938
rect 2168 -5947 2171 -5941
rect 2279 -5939 2283 -5932
rect 2031 -6225 2035 -6081
rect 2052 -6089 2056 -5949
rect 2124 -5957 2202 -5954
rect 2083 -5965 2132 -5961
rect 2083 -5990 2088 -5965
rect 2083 -6045 2088 -5996
rect 2097 -5980 2119 -5975
rect 2097 -5990 2101 -5980
rect 2120 -5990 2124 -5980
rect 2097 -6045 2101 -5996
rect 2106 -6045 2111 -5996
rect 2120 -6045 2124 -5996
rect 2129 -6014 2132 -5965
rect 2142 -5978 2160 -5973
rect 2137 -5990 2142 -5978
rect 2160 -5990 2165 -5978
rect 2129 -6018 2138 -6014
rect 2151 -6023 2155 -5996
rect 2129 -6027 2155 -6023
rect 2106 -6057 2111 -6049
rect 2129 -6057 2132 -6027
rect 2151 -6045 2155 -6027
rect 2174 -6013 2178 -5996
rect 2198 -6012 2202 -5957
rect 2215 -5989 2241 -5984
rect 2217 -5995 2222 -5989
rect 2231 -6012 2235 -6001
rect 2174 -6018 2187 -6013
rect 2198 -6016 2218 -6012
rect 2231 -6016 2265 -6012
rect 2174 -6045 2178 -6018
rect 2231 -6022 2235 -6016
rect 2217 -6035 2221 -6027
rect 2106 -6060 2132 -6057
rect 2209 -6038 2241 -6035
rect 2137 -6060 2141 -6049
rect 2160 -6060 2164 -6049
rect 2137 -6061 2164 -6060
rect 2209 -6061 2212 -6038
rect 2137 -6064 2212 -6061
rect 2148 -6077 2152 -6064
rect 2075 -6080 2152 -6077
rect 2162 -6079 2254 -6076
rect 2172 -6089 2244 -6085
rect 2031 -6387 2035 -6230
rect 2052 -6238 2056 -6094
rect 2123 -6102 2201 -6099
rect 2082 -6110 2131 -6106
rect 2082 -6135 2087 -6110
rect 2064 -6163 2074 -6160
rect 2082 -6190 2087 -6141
rect 2096 -6125 2118 -6120
rect 2096 -6135 2100 -6125
rect 2119 -6135 2123 -6125
rect 2096 -6190 2100 -6141
rect 2105 -6190 2110 -6141
rect 2119 -6190 2123 -6141
rect 2128 -6159 2131 -6110
rect 2141 -6123 2159 -6118
rect 2136 -6135 2141 -6123
rect 2159 -6135 2164 -6123
rect 2128 -6163 2137 -6159
rect 2150 -6168 2154 -6141
rect 2128 -6172 2154 -6168
rect 2105 -6202 2110 -6194
rect 2128 -6202 2131 -6172
rect 2150 -6190 2154 -6172
rect 2173 -6158 2177 -6141
rect 2197 -6157 2201 -6102
rect 2214 -6134 2240 -6129
rect 2216 -6140 2221 -6134
rect 2230 -6157 2234 -6146
rect 2173 -6163 2186 -6158
rect 2197 -6161 2217 -6157
rect 2230 -6161 2251 -6157
rect 2173 -6190 2177 -6163
rect 2230 -6167 2234 -6161
rect 2216 -6180 2220 -6172
rect 2105 -6205 2131 -6202
rect 2208 -6183 2240 -6180
rect 2136 -6205 2140 -6194
rect 2159 -6205 2163 -6194
rect 2136 -6206 2163 -6205
rect 2208 -6206 2211 -6183
rect 2136 -6209 2211 -6206
rect 2147 -6225 2151 -6209
rect 2075 -6228 2151 -6225
rect 2171 -6231 2208 -6228
rect 2233 -6238 2238 -6216
rect 2052 -6242 2238 -6238
rect 2052 -6251 2056 -6242
rect 2148 -6255 2227 -6252
rect 2031 -6539 2035 -6392
rect 2052 -6405 2056 -6256
rect 2123 -6264 2201 -6261
rect 2082 -6272 2131 -6268
rect 2082 -6297 2087 -6272
rect 2064 -6324 2074 -6321
rect 2082 -6352 2087 -6303
rect 2096 -6287 2118 -6282
rect 2096 -6297 2100 -6287
rect 2119 -6297 2123 -6287
rect 2096 -6352 2100 -6303
rect 2105 -6352 2110 -6303
rect 2119 -6352 2123 -6303
rect 2128 -6321 2131 -6272
rect 2141 -6285 2159 -6280
rect 2136 -6297 2141 -6285
rect 2159 -6297 2164 -6285
rect 2128 -6325 2137 -6321
rect 2150 -6330 2154 -6303
rect 2128 -6334 2154 -6330
rect 2105 -6364 2110 -6356
rect 2128 -6364 2131 -6334
rect 2150 -6352 2154 -6334
rect 2173 -6320 2177 -6303
rect 2197 -6319 2201 -6264
rect 2214 -6296 2240 -6291
rect 2216 -6302 2221 -6296
rect 2251 -6301 2256 -6161
rect 2266 -6248 2272 -6016
rect 2279 -6226 2282 -5939
rect 2524 -5943 2529 -5932
rect 2291 -5949 2529 -5943
rect 2291 -6224 2295 -5949
rect 2546 -5958 2549 -5932
rect 2303 -5963 2546 -5959
rect 2303 -6011 2307 -5963
rect 2308 -6016 2499 -6011
rect 2579 -6025 2584 -5930
rect 2579 -6026 2714 -6025
rect 2305 -6032 2714 -6026
rect 2306 -6156 2311 -6032
rect 2759 -6054 2765 -5923
rect 2516 -6060 2765 -6054
rect 2786 -5923 2898 -5917
rect 2311 -6161 2495 -6156
rect 2344 -6216 2495 -6212
rect 2346 -6222 2351 -6216
rect 2369 -6222 2374 -6216
rect 2392 -6222 2397 -6216
rect 2415 -6222 2420 -6216
rect 2471 -6222 2476 -6216
rect 2360 -6238 2364 -6228
rect 2383 -6238 2387 -6228
rect 2406 -6238 2410 -6228
rect 2429 -6238 2433 -6228
rect 2485 -6238 2489 -6228
rect 2360 -6242 2472 -6238
rect 2485 -6242 2495 -6238
rect 2266 -6252 2347 -6248
rect 2429 -6259 2433 -6242
rect 2485 -6259 2489 -6242
rect 2341 -6264 2346 -6259
rect 2364 -6264 2369 -6259
rect 2387 -6264 2392 -6259
rect 2410 -6264 2415 -6259
rect 2341 -6271 2345 -6264
rect 2471 -6273 2475 -6264
rect 2345 -6276 2475 -6273
rect 2376 -6301 2381 -6283
rect 2251 -6307 2381 -6301
rect 2230 -6319 2234 -6308
rect 2400 -6318 2404 -6283
rect 2243 -6319 2400 -6318
rect 2173 -6325 2186 -6320
rect 2197 -6323 2217 -6319
rect 2230 -6323 2400 -6319
rect 2423 -6321 2427 -6284
rect 2173 -6352 2177 -6325
rect 2230 -6329 2234 -6323
rect 2216 -6342 2220 -6334
rect 2105 -6367 2131 -6364
rect 2208 -6345 2240 -6342
rect 2136 -6367 2140 -6356
rect 2159 -6367 2163 -6356
rect 2136 -6368 2163 -6367
rect 2208 -6368 2211 -6345
rect 2136 -6371 2211 -6368
rect 2147 -6385 2151 -6371
rect 2147 -6387 2339 -6385
rect 2075 -6390 2339 -6387
rect 2150 -6399 2361 -6396
rect 2172 -6410 2362 -6407
rect 2031 -6706 2035 -6544
rect 2052 -6645 2056 -6410
rect 2124 -6418 2202 -6415
rect 2083 -6426 2132 -6422
rect 2083 -6451 2088 -6426
rect 2064 -6478 2075 -6474
rect 2083 -6506 2088 -6457
rect 2097 -6441 2119 -6436
rect 2097 -6451 2101 -6441
rect 2120 -6451 2124 -6441
rect 2097 -6506 2101 -6457
rect 2106 -6506 2111 -6457
rect 2120 -6506 2124 -6457
rect 2129 -6475 2132 -6426
rect 2142 -6439 2160 -6434
rect 2137 -6451 2142 -6439
rect 2160 -6451 2165 -6439
rect 2129 -6479 2138 -6475
rect 2151 -6484 2155 -6457
rect 2129 -6488 2155 -6484
rect 2106 -6518 2111 -6510
rect 2129 -6518 2132 -6488
rect 2151 -6506 2155 -6488
rect 2174 -6474 2178 -6457
rect 2198 -6473 2202 -6418
rect 2215 -6450 2241 -6445
rect 2217 -6456 2222 -6450
rect 2231 -6473 2235 -6462
rect 2423 -6472 2428 -6321
rect 2516 -6405 2520 -6060
rect 2786 -6071 2793 -5923
rect 2922 -5958 2925 -5923
rect 2804 -5962 2925 -5958
rect 2944 -6025 2949 -5924
rect 2808 -6032 2949 -6025
rect 2967 -5923 2968 -5918
rect 2529 -6075 2793 -6071
rect 2529 -6394 2533 -6075
rect 2967 -6095 2973 -5923
rect 2542 -6101 2973 -6095
rect 2542 -6102 2971 -6101
rect 2542 -6318 2547 -6102
rect 2596 -6126 2597 -6122
rect 2244 -6473 2429 -6472
rect 2174 -6479 2187 -6474
rect 2198 -6477 2218 -6473
rect 2231 -6477 2429 -6473
rect 2174 -6506 2178 -6479
rect 2231 -6483 2235 -6477
rect 2387 -6478 2429 -6477
rect 2217 -6496 2221 -6488
rect 2106 -6521 2132 -6518
rect 2209 -6499 2241 -6496
rect 2137 -6521 2141 -6510
rect 2160 -6521 2164 -6510
rect 2137 -6522 2164 -6521
rect 2209 -6522 2212 -6499
rect 2137 -6525 2212 -6522
rect 2149 -6541 2153 -6525
rect 2075 -6544 2153 -6541
rect 2596 -6570 2604 -6126
rect 2660 -6156 2666 -6155
rect 2624 -6161 2668 -6156
rect 2402 -6571 2607 -6570
rect 2402 -6574 2642 -6571
rect 2662 -6624 2668 -6161
rect 2683 -6615 2687 -6411
rect 2714 -6571 2720 -6323
rect 2714 -6577 2970 -6571
rect 2702 -6597 2948 -6593
rect 2683 -6619 2895 -6615
rect 2662 -6628 2664 -6624
rect 2670 -6628 2924 -6624
rect 2920 -6637 2924 -6628
rect 2943 -6636 2948 -6597
rect 2965 -6635 2970 -6577
rect 3067 -6640 3196 -6636
rect 3067 -6641 3104 -6640
rect 3067 -6644 3072 -6641
rect 2752 -6645 3072 -6644
rect 2052 -6648 3072 -6645
rect 3099 -6648 3104 -6641
rect 3191 -6648 3196 -6640
rect 2052 -6649 2470 -6648
rect 2081 -6655 2085 -6649
rect 2135 -6655 2140 -6649
rect 2158 -6655 2163 -6649
rect 2214 -6655 2219 -6649
rect 2272 -6654 2277 -6649
rect 2081 -6660 2112 -6655
rect 2088 -6666 2093 -6660
rect 2272 -6659 2303 -6654
rect 2344 -6655 2349 -6649
rect 2367 -6655 2372 -6649
rect 2390 -6655 2395 -6649
rect 2446 -6655 2451 -6649
rect 2499 -6654 2504 -6648
rect 2560 -6649 2756 -6648
rect 2102 -6683 2106 -6672
rect 2149 -6671 2153 -6661
rect 2172 -6671 2176 -6661
rect 2228 -6671 2232 -6661
rect 2279 -6665 2284 -6659
rect 2499 -6659 2530 -6654
rect 2590 -6655 2595 -6649
rect 2613 -6655 2618 -6649
rect 2636 -6655 2641 -6649
rect 2659 -6655 2664 -6649
rect 2715 -6655 2720 -6649
rect 2770 -6654 2774 -6648
rect 2867 -6654 2872 -6648
rect 2890 -6654 2895 -6648
rect 2913 -6654 2918 -6648
rect 2936 -6654 2941 -6648
rect 2959 -6654 2964 -6648
rect 3015 -6654 3020 -6648
rect 3117 -6654 3122 -6648
rect 3140 -6654 3145 -6648
rect 3163 -6654 3168 -6648
rect 2149 -6675 2215 -6671
rect 2228 -6675 2236 -6671
rect 2358 -6670 2362 -6661
rect 2381 -6670 2385 -6661
rect 2404 -6670 2408 -6661
rect 2111 -6683 2136 -6681
rect 2072 -6687 2089 -6683
rect 2102 -6685 2136 -6683
rect 2102 -6687 2115 -6685
rect 2102 -6693 2106 -6687
rect 2172 -6692 2176 -6675
rect 2228 -6692 2232 -6675
rect 2293 -6682 2297 -6671
rect 2304 -6674 2341 -6670
rect 2358 -6671 2408 -6670
rect 2460 -6671 2464 -6661
rect 2506 -6665 2511 -6659
rect 2770 -6659 2801 -6654
rect 2358 -6673 2447 -6671
rect 2304 -6682 2307 -6674
rect 2404 -6675 2447 -6673
rect 2460 -6675 2467 -6671
rect 2604 -6670 2608 -6661
rect 2627 -6670 2631 -6661
rect 2650 -6670 2654 -6661
rect 2673 -6670 2677 -6661
rect 2263 -6686 2280 -6682
rect 2293 -6686 2307 -6682
rect 2310 -6680 2368 -6677
rect 2293 -6692 2297 -6686
rect 2310 -6689 2313 -6680
rect 2153 -6697 2158 -6692
rect 2302 -6692 2313 -6689
rect 2404 -6692 2408 -6675
rect 2460 -6692 2464 -6675
rect 2520 -6682 2524 -6671
rect 2533 -6674 2590 -6670
rect 2604 -6671 2677 -6670
rect 2729 -6671 2733 -6661
rect 2777 -6665 2782 -6659
rect 2604 -6673 2716 -6671
rect 2533 -6682 2537 -6674
rect 2483 -6686 2507 -6682
rect 2520 -6686 2537 -6682
rect 2673 -6675 2716 -6673
rect 2729 -6675 2742 -6671
rect 2520 -6692 2524 -6686
rect 2673 -6692 2677 -6675
rect 2729 -6692 2733 -6675
rect 2791 -6682 2795 -6671
rect 2881 -6670 2885 -6660
rect 2904 -6670 2908 -6660
rect 2927 -6670 2931 -6660
rect 2950 -6670 2954 -6660
rect 2973 -6670 2977 -6660
rect 3029 -6669 3033 -6660
rect 3182 -6666 3186 -6654
rect 3205 -6666 3209 -6654
rect 2881 -6674 3016 -6670
rect 3029 -6673 3093 -6669
rect 3113 -6670 3192 -6666
rect 3205 -6670 3215 -6666
rect 2858 -6682 2868 -6680
rect 2763 -6686 2778 -6682
rect 2791 -6685 2868 -6682
rect 2791 -6686 2859 -6685
rect 2791 -6692 2795 -6686
rect 2973 -6691 2977 -6674
rect 3029 -6691 3033 -6673
rect 3113 -6677 3117 -6670
rect 3136 -6677 3140 -6670
rect 3159 -6677 3163 -6670
rect 3182 -6677 3186 -6670
rect 3205 -6677 3209 -6670
rect 3099 -6689 3103 -6682
rect 3122 -6689 3126 -6682
rect 3145 -6689 3149 -6682
rect 3168 -6689 3172 -6682
rect 3191 -6689 3195 -6682
rect 2302 -6697 2305 -6692
rect 2362 -6697 2367 -6692
rect 2385 -6697 2390 -6692
rect 2608 -6697 2613 -6692
rect 2631 -6697 2636 -6692
rect 2654 -6697 2659 -6692
rect 2885 -6696 2890 -6691
rect 2908 -6696 2913 -6691
rect 2931 -6696 2936 -6691
rect 2954 -6696 2959 -6691
rect 3090 -6693 3195 -6689
rect 2088 -6706 2092 -6698
rect 2135 -6706 2139 -6697
rect 2214 -6706 2218 -6697
rect 2279 -6706 2283 -6697
rect 2344 -6706 2348 -6697
rect 2446 -6706 2450 -6697
rect 2506 -6706 2510 -6697
rect 2590 -6706 2594 -6697
rect 2715 -6706 2719 -6697
rect 2777 -6705 2781 -6697
rect 2867 -6705 2871 -6696
rect 3015 -6704 3019 -6696
rect 3090 -6704 3094 -6693
rect 3015 -6705 3094 -6704
rect 2752 -6706 3094 -6705
rect 2031 -6708 3094 -6706
rect 2031 -6709 2868 -6708
rect 2022 -6724 2066 -6719
rect 2014 -6738 2165 -6733
rect 2257 -6748 2262 -6722
rect 1998 -6753 2262 -6748
rect 2300 -6764 2305 -6721
rect 1986 -6770 2305 -6764
rect 2478 -6789 2483 -6727
rect 1970 -6794 2483 -6789
rect 2764 -6726 2765 -6724
rect 2621 -6802 2625 -6726
rect 2598 -6803 2625 -6802
rect 2412 -6804 2625 -6803
rect 1954 -6807 2625 -6804
rect 2760 -6812 2765 -6726
rect 3129 -6730 3133 -6707
rect 2783 -6735 3133 -6730
rect 3153 -6741 3157 -6707
rect 2784 -6746 3157 -6741
rect 3153 -6747 3157 -6746
rect 3176 -6771 3180 -6703
rect 2790 -6776 3180 -6771
rect 1941 -6816 2765 -6812
<< m2contact >>
rect 517 -4989 523 -4984
rect 609 -5071 618 -5062
rect 720 -5065 726 -5060
rect 775 -5080 781 -5074
rect 922 -5107 927 -5101
rect 958 -5106 963 -5101
rect 1045 -5106 1050 -5101
rect 1148 -5081 1153 -5076
rect 1106 -5089 1111 -5084
rect 1137 -5089 1142 -5084
rect 1238 -5090 1243 -5085
rect 963 -5167 970 -5162
rect 1030 -5167 1035 -5162
rect 1100 -5138 1105 -5133
rect 1169 -5129 1174 -5124
rect 1374 -5090 1379 -5085
rect 1136 -5157 1141 -5152
rect 1052 -5175 1057 -5170
rect 945 -5185 950 -5179
rect 1512 -5090 1517 -5085
rect 1327 -5139 1332 -5134
rect 1158 -5183 1163 -5178
rect 1448 -5183 1453 -5178
rect 1052 -5196 1057 -5191
rect 1790 -5129 1798 -5122
rect 1475 -5183 1480 -5178
rect 1792 -5174 1800 -5167
rect 1100 -5206 1105 -5201
rect 1135 -5206 1140 -5201
rect 1307 -5214 1312 -5209
rect 1169 -5225 1174 -5220
rect 655 -5340 660 -5335
rect -497 -5367 -491 -5362
rect -387 -5367 -381 -5362
rect -275 -5366 -269 -5361
rect -163 -5366 -157 -5361
rect -52 -5366 -46 -5361
rect 60 -5367 66 -5362
rect 172 -5367 178 -5362
rect 764 -5341 769 -5334
rect 875 -5341 880 -5335
rect 986 -5342 992 -5336
rect 1099 -5340 1104 -5335
rect 1211 -5341 1216 -5336
rect 1323 -5341 1328 -5336
rect 1435 -5341 1442 -5334
rect 1875 -5338 1881 -5333
rect 1983 -5339 1989 -5334
rect 2095 -5339 2101 -5334
rect 2208 -5339 2214 -5334
rect 2318 -5339 2324 -5334
rect 2429 -5339 2435 -5334
rect 2542 -5339 2548 -5334
rect 2655 -5339 2661 -5334
rect 283 -5367 289 -5362
rect 2668 -5372 2674 -5367
rect 1260 -5602 1272 -5593
rect -623 -5785 -618 -5780
rect -497 -5613 -490 -5608
rect -388 -5610 -381 -5605
rect -521 -5637 -514 -5631
rect -276 -5612 -269 -5607
rect -381 -5661 -372 -5654
rect -164 -5613 -157 -5608
rect -244 -5686 -236 -5677
rect 514 -5635 526 -5623
rect 926 -5665 936 -5652
rect 596 -5679 605 -5673
rect 703 -5677 714 -5668
rect 814 -5675 825 -5667
rect -95 -5705 -87 -5697
rect -1880 -5866 -1871 -5857
rect -623 -5813 -618 -5808
rect -1787 -5866 -1778 -5857
rect 1376 -5605 1386 -5599
rect 1328 -6015 1345 -5998
rect 1778 -5619 1788 -5608
rect 1376 -6047 1388 -6035
rect -1880 -6281 -1869 -6271
rect -1569 -6267 -1564 -6262
rect -1796 -6280 -1785 -6270
rect -779 -6267 -773 -6262
rect 202 -6267 209 -6262
rect 1087 -6266 1093 -6261
rect -779 -6287 -773 -6282
rect 203 -6286 210 -6281
rect -1569 -6295 -1564 -6290
rect -1509 -6308 -1501 -6300
rect -711 -6307 -697 -6297
rect 142 -6300 150 -6293
rect 1086 -6290 1095 -6283
rect 1020 -6309 1027 -6302
rect -1603 -6508 -1598 -6503
rect -1787 -6613 -1782 -6608
rect -1617 -6575 -1612 -6570
rect -1533 -6469 -1528 -6464
rect -1414 -6454 -1409 -6449
rect -1525 -6508 -1520 -6503
rect -1575 -6575 -1570 -6570
rect -1485 -6564 -1480 -6559
rect -1555 -6584 -1550 -6579
rect -1485 -6602 -1480 -6597
rect -1651 -6613 -1646 -6608
rect -1698 -6640 -1693 -6635
rect -1698 -6661 -1693 -6656
rect -1614 -6686 -1609 -6681
rect -1555 -6610 -1550 -6605
rect -1520 -6613 -1515 -6608
rect -1536 -6686 -1531 -6681
rect -1474 -6684 -1469 -6679
rect -1378 -6613 -1373 -6608
rect -1391 -6683 -1386 -6678
rect -802 -6506 -797 -6501
rect -986 -6611 -981 -6606
rect -816 -6573 -811 -6568
rect -732 -6467 -727 -6462
rect -613 -6452 -608 -6447
rect -724 -6506 -719 -6501
rect -774 -6573 -769 -6568
rect -684 -6562 -679 -6557
rect -754 -6582 -749 -6577
rect -684 -6600 -679 -6595
rect -850 -6611 -845 -6606
rect -897 -6638 -892 -6633
rect -897 -6659 -892 -6654
rect -964 -6685 -953 -6675
rect -813 -6684 -808 -6679
rect -754 -6608 -749 -6603
rect -719 -6611 -714 -6606
rect -735 -6684 -730 -6679
rect -673 -6682 -668 -6677
rect -577 -6611 -572 -6606
rect -590 -6681 -585 -6676
rect 101 -6506 106 -6501
rect -83 -6611 -78 -6606
rect 87 -6573 92 -6568
rect 171 -6467 176 -6462
rect 290 -6452 295 -6447
rect 179 -6506 184 -6501
rect 129 -6573 134 -6568
rect 219 -6562 224 -6557
rect 149 -6582 154 -6577
rect 219 -6600 224 -6595
rect 53 -6611 58 -6606
rect 6 -6638 11 -6633
rect 6 -6659 11 -6654
rect -60 -6688 -49 -6678
rect 90 -6684 95 -6679
rect 149 -6608 154 -6603
rect 184 -6611 189 -6606
rect 168 -6684 173 -6679
rect 230 -6682 235 -6677
rect 326 -6611 331 -6606
rect 313 -6681 318 -6676
rect 969 -6505 974 -6500
rect 785 -6610 790 -6605
rect 955 -6572 960 -6567
rect 1039 -6466 1044 -6461
rect 1158 -6451 1163 -6446
rect 1047 -6505 1052 -6500
rect 2094 -5603 2103 -5593
rect 1833 -5619 1843 -5608
rect 2206 -5616 2218 -5606
rect 2733 -5372 2740 -5367
rect 1872 -5756 1884 -5747
rect 1982 -5775 1990 -5768
rect 2031 -5754 2036 -5749
rect 2100 -5754 2105 -5749
rect 2170 -5774 2179 -5768
rect 2899 -5772 2904 -5767
rect 2370 -5785 2378 -5780
rect 2245 -5830 2250 -5825
rect 2543 -5800 2548 -5793
rect 2469 -5831 2474 -5826
rect 2741 -5834 2746 -5829
rect 2032 -5902 2037 -5897
rect 2014 -5936 2019 -5931
rect 1986 -6164 1991 -6159
rect 1954 -6325 1959 -6320
rect 1915 -6479 1926 -6471
rect 997 -6572 1002 -6567
rect 1087 -6561 1092 -6556
rect 1017 -6581 1022 -6576
rect 1087 -6599 1092 -6594
rect 921 -6610 926 -6605
rect 874 -6637 879 -6632
rect 874 -6658 879 -6653
rect 809 -6687 819 -6678
rect 958 -6683 963 -6678
rect 1017 -6607 1022 -6602
rect 1052 -6610 1057 -6605
rect 1036 -6683 1041 -6678
rect 1098 -6681 1103 -6676
rect 1194 -6610 1199 -6605
rect 1181 -6680 1186 -6675
rect -964 -6813 -953 -6803
rect -60 -6813 -49 -6803
rect 809 -6813 820 -6803
rect 2022 -5910 2027 -5905
rect 2031 -6081 2036 -6076
rect 2244 -5867 2249 -5862
rect 2468 -5867 2473 -5862
rect 2245 -5879 2250 -5874
rect 2086 -5902 2091 -5897
rect 2299 -5894 2304 -5889
rect 2309 -5894 2314 -5889
rect 2741 -5867 2746 -5862
rect 2472 -5879 2477 -5874
rect 2759 -5880 2765 -5875
rect 2528 -5895 2533 -5890
rect 2545 -5895 2550 -5890
rect 2106 -5909 2111 -5904
rect 2065 -5936 2070 -5931
rect 2471 -5932 2476 -5927
rect 2524 -5932 2529 -5927
rect 2545 -5932 2550 -5927
rect 2759 -5923 2765 -5918
rect 2052 -5949 2057 -5944
rect 2119 -5958 2124 -5953
rect 2119 -5980 2124 -5975
rect 2137 -5978 2142 -5973
rect 2160 -5978 2165 -5973
rect 2210 -5989 2215 -5984
rect 2265 -6016 2272 -6011
rect 2070 -6081 2075 -6076
rect 2254 -6079 2259 -6074
rect 2052 -6094 2057 -6089
rect 2244 -6090 2249 -6085
rect 2031 -6230 2036 -6225
rect 2118 -6103 2123 -6098
rect 2059 -6164 2064 -6159
rect 2118 -6125 2123 -6120
rect 2136 -6123 2141 -6118
rect 2159 -6123 2164 -6118
rect 2209 -6134 2214 -6129
rect 2251 -6161 2256 -6156
rect 2070 -6230 2075 -6225
rect 2233 -6216 2238 -6211
rect 2208 -6231 2213 -6226
rect 2052 -6256 2057 -6251
rect 2227 -6256 2232 -6251
rect 2031 -6392 2036 -6387
rect 2118 -6265 2123 -6260
rect 2059 -6325 2064 -6320
rect 2118 -6287 2123 -6282
rect 2136 -6285 2141 -6280
rect 2159 -6285 2164 -6280
rect 2209 -6296 2214 -6291
rect 2546 -5963 2551 -5958
rect 2301 -6016 2308 -6011
rect 2499 -6016 2504 -6011
rect 2714 -6032 2723 -6025
rect 2306 -6161 2311 -6156
rect 2495 -6161 2500 -6156
rect 2339 -6216 2344 -6211
rect 2278 -6231 2283 -6226
rect 2291 -6229 2296 -6224
rect 2340 -6276 2345 -6271
rect 2400 -6323 2405 -6318
rect 2070 -6392 2075 -6387
rect 2339 -6390 2344 -6385
rect 2361 -6399 2366 -6394
rect 2052 -6410 2057 -6405
rect 2362 -6410 2367 -6405
rect 2031 -6544 2036 -6539
rect 2119 -6419 2124 -6414
rect 2059 -6478 2064 -6473
rect 2119 -6441 2124 -6436
rect 2137 -6439 2142 -6434
rect 2160 -6439 2165 -6434
rect 2210 -6450 2215 -6445
rect 2798 -5962 2804 -5957
rect 2803 -6032 2808 -6025
rect 2542 -6323 2547 -6318
rect 2597 -6126 2606 -6119
rect 2528 -6399 2533 -6394
rect 2515 -6410 2520 -6405
rect 2070 -6544 2075 -6539
rect 2618 -6161 2624 -6156
rect 2713 -6323 2721 -6318
rect 2683 -6411 2688 -6406
rect 2236 -6675 2242 -6670
rect 2067 -6688 2072 -6683
rect 2467 -6675 2472 -6670
rect 2257 -6687 2263 -6682
rect 2478 -6686 2483 -6681
rect 2742 -6675 2747 -6670
rect 2757 -6687 2763 -6682
rect 2301 -6702 2306 -6697
rect 2066 -6724 2071 -6719
rect 2257 -6722 2262 -6717
rect 2300 -6721 2305 -6716
rect 2478 -6727 2483 -6722
rect 2758 -6726 2764 -6721
rect 2777 -6735 2783 -6730
rect 2778 -6746 2784 -6741
rect 2784 -6776 2790 -6771
<< metal2 >>
rect -495 -5608 -492 -5367
rect -386 -5605 -383 -5367
rect -274 -5607 -271 -5366
rect -162 -5608 -159 -5366
rect -51 -5632 -48 -5366
rect -514 -5636 -48 -5632
rect 61 -5656 64 -5367
rect -372 -5660 65 -5656
rect 173 -5679 176 -5367
rect -236 -5685 177 -5679
rect 285 -5697 288 -5367
rect 517 -5623 523 -4989
rect 610 -5179 617 -5071
rect 720 -5162 726 -5065
rect 781 -5079 1148 -5076
rect 1047 -5088 1106 -5085
rect 1047 -5101 1050 -5088
rect 1142 -5088 1238 -5085
rect 927 -5106 958 -5101
rect 720 -5166 963 -5162
rect 1100 -5163 1103 -5138
rect 1138 -5152 1141 -5089
rect 1243 -5088 1374 -5085
rect 1379 -5088 1512 -5085
rect 1517 -5088 1518 -5085
rect 1035 -5166 1103 -5163
rect 610 -5185 945 -5179
rect 1052 -5191 1057 -5175
rect 1100 -5201 1103 -5166
rect 1158 -5203 1161 -5183
rect 1140 -5206 1161 -5203
rect 1169 -5220 1174 -5129
rect 1307 -5138 1327 -5134
rect 1307 -5209 1310 -5138
rect 1792 -5167 1796 -5129
rect 1453 -5182 1475 -5179
rect 656 -5379 659 -5340
rect 598 -5384 659 -5379
rect 598 -5673 602 -5384
rect 764 -5385 769 -5341
rect 876 -5385 880 -5341
rect 705 -5391 769 -5385
rect 705 -5668 711 -5391
rect 815 -5392 880 -5385
rect 987 -5388 992 -5342
rect 1099 -5386 1103 -5340
rect 1211 -5385 1216 -5341
rect 815 -5667 823 -5392
rect 928 -5395 992 -5388
rect 1002 -5393 1103 -5386
rect 1110 -5392 1216 -5385
rect 1323 -5390 1328 -5341
rect 1436 -5389 1440 -5341
rect 928 -5652 935 -5395
rect -87 -5703 288 -5697
rect -623 -5808 -618 -5785
rect -1871 -5865 -1787 -5859
rect 1002 -5930 1011 -5393
rect -1463 -5939 1011 -5930
rect 1110 -5592 1118 -5392
rect 1261 -5397 1328 -5390
rect 1377 -5394 1440 -5389
rect -1869 -6280 -1796 -6272
rect -1869 -6281 -1785 -6280
rect -1569 -6290 -1564 -6267
rect -1463 -6300 -1455 -5939
rect 1110 -5959 1119 -5592
rect 1261 -5593 1269 -5397
rect 1377 -5599 1384 -5394
rect 1788 -5618 1833 -5608
rect 1876 -5747 1881 -5338
rect 1984 -5768 1989 -5339
rect 2096 -5593 2101 -5339
rect 2208 -5606 2213 -5339
rect 2319 -5643 2324 -5339
rect 2430 -5598 2435 -5339
rect 2172 -5647 2324 -5643
rect 2373 -5602 2435 -5598
rect 2036 -5753 2100 -5750
rect 2172 -5768 2175 -5647
rect 2373 -5780 2376 -5602
rect 2543 -5793 2548 -5339
rect 2655 -5600 2660 -5339
rect 2674 -5372 2733 -5367
rect 2655 -5604 2903 -5600
rect 2900 -5767 2903 -5604
rect 2245 -5862 2248 -5830
rect 2469 -5862 2472 -5831
rect 2742 -5862 2745 -5834
rect 2037 -5901 2086 -5898
rect 2027 -5909 2106 -5906
rect 2019 -5935 2065 -5931
rect 2057 -5949 2141 -5944
rect -658 -5970 1119 -5959
rect -779 -6282 -774 -6267
rect -1501 -6308 -1455 -6300
rect -658 -6298 -651 -5970
rect 2120 -5975 2123 -5958
rect 2137 -5973 2141 -5949
rect 2165 -5977 2214 -5974
rect 2211 -5984 2214 -5977
rect -697 -6306 -651 -6298
rect 142 -6014 1328 -6002
rect 142 -6293 149 -6014
rect 1020 -6044 1376 -6037
rect 204 -6281 208 -6267
rect 1020 -6302 1027 -6044
rect 2036 -6081 2070 -6077
rect 2245 -6085 2249 -5879
rect 2299 -5906 2302 -5894
rect 2254 -5909 2302 -5906
rect 2254 -6074 2258 -5909
rect 2309 -5915 2313 -5894
rect 2266 -5921 2313 -5915
rect 2266 -6011 2272 -5921
rect 2472 -5927 2475 -5879
rect 2524 -5927 2528 -5892
rect 2545 -5927 2549 -5895
rect 2760 -5918 2763 -5880
rect 2551 -5962 2798 -5958
rect 2272 -6016 2301 -6012
rect 2504 -6016 2603 -6011
rect 2057 -6094 2141 -6089
rect 2119 -6120 2122 -6103
rect 2137 -6118 2141 -6094
rect 2597 -6119 2603 -6016
rect 2723 -6032 2803 -6025
rect 2164 -6122 2213 -6119
rect 2210 -6129 2213 -6122
rect 1991 -6163 2059 -6160
rect 2256 -6161 2306 -6156
rect 2500 -6161 2618 -6156
rect 2238 -6215 2339 -6211
rect 2036 -6230 2070 -6226
rect 2213 -6231 2278 -6228
rect 2057 -6256 2140 -6251
rect 2291 -6252 2296 -6229
rect 2232 -6255 2296 -6252
rect 1088 -6283 1092 -6266
rect 2119 -6282 2122 -6265
rect 2136 -6280 2140 -6256
rect 2164 -6284 2213 -6281
rect 2210 -6291 2213 -6284
rect 1959 -6325 2059 -6321
rect 2340 -6385 2344 -6276
rect 2405 -6323 2542 -6318
rect 2547 -6323 2713 -6318
rect 2036 -6392 2070 -6388
rect 2366 -6399 2528 -6395
rect 2057 -6410 2142 -6405
rect 2367 -6410 2515 -6406
rect 2520 -6410 2683 -6406
rect 2120 -6436 2123 -6419
rect 2138 -6434 2142 -6410
rect 2165 -6438 2214 -6435
rect 2211 -6445 2214 -6438
rect -1453 -6453 -1414 -6449
rect -1453 -6456 -1450 -6453
rect -652 -6451 -613 -6447
rect -652 -6454 -649 -6451
rect 251 -6451 290 -6447
rect 251 -6454 254 -6451
rect 1119 -6450 1158 -6446
rect 1119 -6453 1122 -6450
rect -1532 -6460 -1450 -6456
rect -731 -6458 -649 -6454
rect 172 -6458 254 -6454
rect 1040 -6457 1122 -6453
rect -1532 -6464 -1529 -6460
rect -731 -6462 -728 -6458
rect 172 -6462 175 -6458
rect 1040 -6461 1043 -6457
rect 1926 -6478 2059 -6473
rect -1598 -6507 -1525 -6504
rect -797 -6505 -724 -6502
rect 106 -6505 179 -6502
rect 974 -6504 1047 -6501
rect 2036 -6544 2070 -6540
rect -1612 -6574 -1575 -6571
rect -1554 -6605 -1551 -6584
rect -1484 -6597 -1481 -6564
rect -811 -6572 -774 -6569
rect -753 -6603 -750 -6582
rect -683 -6595 -680 -6562
rect 92 -6572 129 -6569
rect 150 -6603 153 -6582
rect 220 -6595 223 -6562
rect 960 -6571 997 -6568
rect 1018 -6602 1021 -6581
rect 1088 -6594 1091 -6561
rect -1782 -6612 -1651 -6609
rect -1646 -6612 -1565 -6609
rect -1568 -6615 -1565 -6612
rect -1541 -6612 -1520 -6609
rect -1541 -6615 -1538 -6612
rect -1515 -6612 -1378 -6609
rect -981 -6610 -850 -6607
rect -845 -6610 -764 -6607
rect -767 -6613 -764 -6610
rect -740 -6610 -719 -6607
rect -740 -6613 -737 -6610
rect -714 -6610 -577 -6607
rect -78 -6610 53 -6607
rect 58 -6610 139 -6607
rect -1568 -6618 -1538 -6615
rect -767 -6616 -737 -6613
rect 136 -6613 139 -6610
rect 163 -6610 184 -6607
rect 163 -6613 166 -6610
rect 189 -6610 326 -6607
rect 790 -6609 921 -6606
rect 926 -6609 1007 -6606
rect 136 -6616 166 -6613
rect 1004 -6612 1007 -6609
rect 1031 -6609 1052 -6606
rect 1031 -6612 1034 -6609
rect 1057 -6609 1194 -6606
rect 1004 -6615 1034 -6612
rect -1697 -6656 -1694 -6640
rect -896 -6654 -893 -6638
rect 7 -6654 10 -6638
rect 875 -6653 878 -6637
rect -1609 -6685 -1536 -6682
rect -1469 -6683 -1391 -6680
rect -808 -6683 -735 -6680
rect -668 -6681 -590 -6678
rect -964 -6803 -954 -6685
rect 95 -6683 168 -6680
rect 235 -6681 313 -6678
rect 963 -6682 1036 -6679
rect 1103 -6680 1181 -6677
rect -60 -6803 -50 -6688
rect 809 -6803 819 -6687
rect 2067 -6719 2071 -6688
rect 2237 -6772 2240 -6675
rect 2257 -6717 2262 -6687
rect 2301 -6716 2304 -6702
rect 2468 -6737 2471 -6675
rect 2478 -6722 2482 -6686
rect 2743 -6731 2746 -6675
rect 2758 -6721 2761 -6687
rect 2743 -6735 2777 -6731
rect 2468 -6740 2666 -6737
rect 2662 -6743 2666 -6740
rect 2662 -6746 2778 -6743
rect 2237 -6776 2784 -6772
<< labels >>
rlabel metal1 1122 -5088 1125 -5086 1 vdd
rlabel metal1 1119 -5206 1123 -5204 1 gnd
rlabel metal1 1044 -5131 1048 -5129 1 D3
rlabel metal1 1570 -5127 1574 -5125 7 D2
rlabel metal1 1414 -5127 1418 -5125 1 D1
rlabel metal1 1282 -5127 1286 -5125 1 D0
rlabel metal1 1105 -5183 1109 -5181 1 S0
rlabel metal1 1106 -5115 1110 -5113 1 S1
rlabel polysilicon -553 -5353 -550 -5350 1 B3
rlabel polysilicon -445 -5352 -442 -5349 1 B2
rlabel polysilicon -333 -5352 -330 -5349 1 B1
rlabel polysilicon -221 -5352 -218 -5349 1 B0
rlabel polysilicon -110 -5351 -107 -5348 1 A3
rlabel polysilicon 2 -5352 5 -5349 1 A2
rlabel polysilicon 114 -5351 117 -5348 1 A1
rlabel polysilicon 226 -5351 229 -5348 1 A0
rlabel metal1 280 -5346 283 -5343 7 A0_out
rlabel metal1 167 -5346 170 -5343 1 A1_out
rlabel metal1 56 -5347 59 -5344 1 A2_out
rlabel metal1 -57 -5347 -54 -5344 1 A3_out
rlabel metal1 -167 -5347 -164 -5344 1 B0_out
rlabel metal1 -279 -5347 -276 -5344 1 B1_out
rlabel metal1 -391 -5347 -388 -5344 1 B2_out
rlabel metal1 -499 -5347 -496 -5344 1 B3_out
rlabel metal1 -42 -5830 -39 -5828 7 Y0
rlabel metal1 -192 -5830 -189 -5828 1 Y1
rlabel metal1 -331 -5830 -328 -5828 1 Y2
rlabel metal1 -469 -5830 -466 -5828 1 Y3
rlabel metal1 2681 -5730 2684 -5728 1 AB
rlabel metal1 2491 -6241 2494 -6239 1 AequalB
rlabel metal1 3211 -6669 3214 -6667 7 BA
rlabel metal1 -1141 -6652 -1138 -6650 7 carry
rlabel metal1 -1391 -6467 -1387 -6465 1 YS3
rlabel metal1 -589 -6465 -586 -6463 1 YS2
rlabel metal1 313 -6464 317 -6463 1 YS1
rlabel metal1 1182 -6463 1185 -6462 1 YS0
rlabel metal1 735 -4989 741 -4986 5 M
rlabel metal1 634 -5032 638 -5030 1 add1
<< end >>
