magic
tech scmos
timestamp 1700160321
<< nwell >>
rect 498 480 621 498
rect 23 331 54 349
rect 70 342 124 360
rect 149 342 180 360
rect 206 332 237 350
rect 271 342 348 360
rect 373 342 404 360
rect 434 332 465 350
rect 518 342 618 360
rect 643 342 674 360
rect 708 331 739 349
rect 798 342 921 360
rect 946 342 977 360
rect 12 199 120 217
rect 146 194 177 212
rect 11 54 119 72
rect 145 49 176 67
rect 275 -33 375 -15
rect 400 -33 431 -15
rect 11 -108 119 -90
rect 145 -113 176 -95
rect 12 -262 120 -244
rect 146 -267 177 -249
rect 17 -477 48 -459
rect 64 -466 118 -448
rect 143 -466 174 -448
rect 208 -476 239 -458
rect 273 -466 350 -448
rect 375 -466 406 -448
rect 435 -476 466 -458
rect 519 -466 619 -448
rect 644 -466 675 -448
rect 706 -476 737 -458
rect 796 -465 919 -447
rect 944 -465 975 -447
rect 1028 -459 1151 -441
<< ntransistor >>
rect 513 458 516 463
rect 536 458 539 463
rect 559 458 562 463
rect 582 458 585 463
rect 605 458 608 463
rect 38 311 41 316
rect 85 312 88 317
rect 108 312 111 317
rect 164 312 167 317
rect 221 312 224 317
rect 286 312 289 317
rect 309 312 312 317
rect 332 312 335 317
rect 388 312 391 317
rect 449 312 452 317
rect 533 312 536 317
rect 556 312 559 317
rect 579 312 582 317
rect 602 312 605 317
rect 658 312 661 317
rect 723 311 726 316
rect 813 312 816 317
rect 836 312 839 317
rect 859 312 862 317
rect 882 312 885 317
rect 905 312 908 317
rect 961 312 964 317
rect 27 152 30 156
rect 50 152 53 156
rect 81 152 84 156
rect 104 152 107 156
rect 161 174 164 179
rect 26 7 29 11
rect 49 7 52 11
rect 80 7 83 11
rect 103 7 106 11
rect 160 29 163 34
rect 290 -63 293 -58
rect 313 -63 316 -58
rect 336 -63 339 -58
rect 359 -63 362 -58
rect 415 -63 418 -58
rect 26 -155 29 -151
rect 49 -155 52 -151
rect 80 -155 83 -151
rect 103 -155 106 -151
rect 160 -133 163 -128
rect 27 -309 30 -305
rect 50 -309 53 -305
rect 81 -309 84 -305
rect 104 -309 107 -305
rect 161 -287 164 -282
rect 1043 -481 1046 -476
rect 1066 -481 1069 -476
rect 1089 -481 1092 -476
rect 1112 -481 1115 -476
rect 1135 -481 1138 -476
rect 32 -497 35 -492
rect 79 -496 82 -491
rect 102 -496 105 -491
rect 158 -496 161 -491
rect 223 -496 226 -491
rect 288 -496 291 -491
rect 311 -496 314 -491
rect 334 -496 337 -491
rect 390 -496 393 -491
rect 450 -496 453 -491
rect 534 -496 537 -491
rect 557 -496 560 -491
rect 580 -496 583 -491
rect 603 -496 606 -491
rect 659 -496 662 -491
rect 721 -496 724 -491
rect 811 -495 814 -490
rect 834 -495 837 -490
rect 857 -495 860 -490
rect 880 -495 883 -490
rect 903 -495 906 -490
rect 959 -495 962 -490
<< ptransistor >>
rect 513 486 516 492
rect 536 486 539 492
rect 559 486 562 492
rect 582 486 585 492
rect 605 486 608 492
rect 85 348 88 354
rect 108 348 111 354
rect 164 348 167 354
rect 286 348 289 354
rect 309 348 312 354
rect 332 348 335 354
rect 388 348 391 354
rect 533 348 536 354
rect 556 348 559 354
rect 579 348 582 354
rect 602 348 605 354
rect 658 348 661 354
rect 813 348 816 354
rect 836 348 839 354
rect 859 348 862 354
rect 882 348 885 354
rect 905 348 908 354
rect 961 348 964 354
rect 38 337 41 343
rect 221 338 224 344
rect 449 338 452 344
rect 723 337 726 343
rect 27 205 30 211
rect 50 205 53 211
rect 81 205 84 211
rect 104 205 107 211
rect 161 200 164 206
rect 26 60 29 66
rect 49 60 52 66
rect 80 60 83 66
rect 103 60 106 66
rect 160 55 163 61
rect 290 -27 293 -21
rect 313 -27 316 -21
rect 336 -27 339 -21
rect 359 -27 362 -21
rect 415 -27 418 -21
rect 26 -102 29 -96
rect 49 -102 52 -96
rect 80 -102 83 -96
rect 103 -102 106 -96
rect 160 -107 163 -101
rect 27 -256 30 -250
rect 50 -256 53 -250
rect 81 -256 84 -250
rect 104 -256 107 -250
rect 161 -261 164 -255
rect 1043 -453 1046 -447
rect 1066 -453 1069 -447
rect 1089 -453 1092 -447
rect 1112 -453 1115 -447
rect 1135 -453 1138 -447
rect 79 -460 82 -454
rect 102 -460 105 -454
rect 158 -460 161 -454
rect 288 -460 291 -454
rect 311 -460 314 -454
rect 334 -460 337 -454
rect 390 -460 393 -454
rect 534 -460 537 -454
rect 557 -460 560 -454
rect 580 -460 583 -454
rect 603 -460 606 -454
rect 659 -460 662 -454
rect 811 -459 814 -453
rect 834 -459 837 -453
rect 857 -459 860 -453
rect 880 -459 883 -453
rect 903 -459 906 -453
rect 959 -459 962 -453
rect 32 -471 35 -465
rect 223 -470 226 -464
rect 450 -470 453 -464
rect 721 -470 724 -464
<< ndiffusion >>
rect 509 458 513 463
rect 516 458 519 463
rect 532 458 536 463
rect 539 458 542 463
rect 555 458 559 463
rect 562 458 565 463
rect 578 458 582 463
rect 585 458 588 463
rect 601 458 605 463
rect 608 458 611 463
rect 34 311 38 316
rect 41 311 44 316
rect 81 312 85 317
rect 88 312 91 317
rect 104 312 108 317
rect 111 312 114 317
rect 160 312 164 317
rect 167 312 170 317
rect 217 312 221 317
rect 224 312 227 317
rect 282 312 286 317
rect 289 312 292 317
rect 305 312 309 317
rect 312 312 315 317
rect 328 312 332 317
rect 335 312 338 317
rect 384 312 388 317
rect 391 312 394 317
rect 445 312 449 317
rect 452 312 455 317
rect 529 312 533 317
rect 536 312 539 317
rect 552 312 556 317
rect 559 312 562 317
rect 575 312 579 317
rect 582 312 585 317
rect 598 312 602 317
rect 605 312 608 317
rect 654 312 658 317
rect 661 312 664 317
rect 719 311 723 316
rect 726 311 729 316
rect 809 312 813 317
rect 816 312 819 317
rect 832 312 836 317
rect 839 312 842 317
rect 855 312 859 317
rect 862 312 865 317
rect 878 312 882 317
rect 885 312 888 317
rect 901 312 905 317
rect 908 312 911 317
rect 957 312 961 317
rect 964 312 967 317
rect 24 152 27 156
rect 30 152 33 156
rect 47 152 50 156
rect 53 152 56 156
rect 77 152 81 156
rect 84 152 87 156
rect 100 152 104 156
rect 107 152 110 156
rect 157 174 161 179
rect 164 174 167 179
rect 23 7 26 11
rect 29 7 32 11
rect 46 7 49 11
rect 52 7 55 11
rect 76 7 80 11
rect 83 7 86 11
rect 99 7 103 11
rect 106 7 109 11
rect 156 29 160 34
rect 163 29 166 34
rect 286 -63 290 -58
rect 293 -63 296 -58
rect 309 -63 313 -58
rect 316 -63 319 -58
rect 332 -63 336 -58
rect 339 -63 342 -58
rect 355 -63 359 -58
rect 362 -63 365 -58
rect 411 -63 415 -58
rect 418 -63 421 -58
rect 23 -155 26 -151
rect 29 -155 32 -151
rect 46 -155 49 -151
rect 52 -155 55 -151
rect 76 -155 80 -151
rect 83 -155 86 -151
rect 99 -155 103 -151
rect 106 -155 109 -151
rect 156 -133 160 -128
rect 163 -133 166 -128
rect 24 -309 27 -305
rect 30 -309 33 -305
rect 47 -309 50 -305
rect 53 -309 56 -305
rect 77 -309 81 -305
rect 84 -309 87 -305
rect 100 -309 104 -305
rect 107 -309 110 -305
rect 157 -287 161 -282
rect 164 -287 167 -282
rect 1039 -481 1043 -476
rect 1046 -481 1049 -476
rect 1062 -481 1066 -476
rect 1069 -481 1072 -476
rect 1085 -481 1089 -476
rect 1092 -481 1095 -476
rect 1108 -481 1112 -476
rect 1115 -481 1118 -476
rect 1131 -481 1135 -476
rect 1138 -481 1141 -476
rect 28 -497 32 -492
rect 35 -497 38 -492
rect 75 -496 79 -491
rect 82 -496 85 -491
rect 98 -496 102 -491
rect 105 -496 108 -491
rect 154 -496 158 -491
rect 161 -496 164 -491
rect 219 -496 223 -491
rect 226 -496 229 -491
rect 284 -496 288 -491
rect 291 -496 294 -491
rect 307 -496 311 -491
rect 314 -496 317 -491
rect 330 -496 334 -491
rect 337 -496 340 -491
rect 386 -496 390 -491
rect 393 -496 396 -491
rect 446 -496 450 -491
rect 453 -496 456 -491
rect 530 -496 534 -491
rect 537 -496 540 -491
rect 553 -496 557 -491
rect 560 -496 563 -491
rect 576 -496 580 -491
rect 583 -496 586 -491
rect 599 -496 603 -491
rect 606 -496 609 -491
rect 655 -496 659 -491
rect 662 -496 665 -491
rect 717 -496 721 -491
rect 724 -496 727 -491
rect 807 -495 811 -490
rect 814 -495 817 -490
rect 830 -495 834 -490
rect 837 -495 840 -490
rect 853 -495 857 -490
rect 860 -495 863 -490
rect 876 -495 880 -490
rect 883 -495 886 -490
rect 899 -495 903 -490
rect 906 -495 909 -490
rect 955 -495 959 -490
rect 962 -495 965 -490
<< pdiffusion >>
rect 510 486 513 492
rect 516 486 519 492
rect 533 486 536 492
rect 539 486 542 492
rect 556 486 559 492
rect 562 486 565 492
rect 579 486 582 492
rect 585 486 588 492
rect 602 486 605 492
rect 608 486 611 492
rect 82 348 85 354
rect 88 348 91 354
rect 105 348 108 354
rect 111 348 114 354
rect 161 348 164 354
rect 167 348 170 354
rect 283 348 286 354
rect 289 348 292 354
rect 306 348 309 354
rect 312 348 315 354
rect 329 348 332 354
rect 335 348 338 354
rect 385 348 388 354
rect 391 348 394 354
rect 530 348 533 354
rect 536 348 539 354
rect 553 348 556 354
rect 559 348 562 354
rect 576 348 579 354
rect 582 348 585 354
rect 599 348 602 354
rect 605 348 608 354
rect 655 348 658 354
rect 661 348 664 354
rect 810 348 813 354
rect 816 348 819 354
rect 833 348 836 354
rect 839 348 842 354
rect 856 348 859 354
rect 862 348 865 354
rect 879 348 882 354
rect 885 348 888 354
rect 902 348 905 354
rect 908 348 911 354
rect 958 348 961 354
rect 964 348 967 354
rect 35 337 38 343
rect 41 337 44 343
rect 218 338 221 344
rect 224 338 227 344
rect 446 338 449 344
rect 452 338 455 344
rect 720 337 723 343
rect 726 337 729 343
rect 24 205 27 211
rect 30 205 33 211
rect 47 205 50 211
rect 53 205 56 211
rect 78 205 81 211
rect 84 205 87 211
rect 101 205 104 211
rect 107 205 110 211
rect 158 200 161 206
rect 164 200 167 206
rect 23 60 26 66
rect 29 60 32 66
rect 46 60 49 66
rect 52 60 55 66
rect 77 60 80 66
rect 83 60 86 66
rect 100 60 103 66
rect 106 60 109 66
rect 157 55 160 61
rect 163 55 166 61
rect 287 -27 290 -21
rect 293 -27 296 -21
rect 310 -27 313 -21
rect 316 -27 319 -21
rect 333 -27 336 -21
rect 339 -27 342 -21
rect 356 -27 359 -21
rect 362 -27 365 -21
rect 412 -27 415 -21
rect 418 -27 421 -21
rect 23 -102 26 -96
rect 29 -102 32 -96
rect 46 -102 49 -96
rect 52 -102 55 -96
rect 77 -102 80 -96
rect 83 -102 86 -96
rect 100 -102 103 -96
rect 106 -102 109 -96
rect 157 -107 160 -101
rect 163 -107 166 -101
rect 24 -256 27 -250
rect 30 -256 33 -250
rect 47 -256 50 -250
rect 53 -256 56 -250
rect 78 -256 81 -250
rect 84 -256 87 -250
rect 101 -256 104 -250
rect 107 -256 110 -250
rect 158 -261 161 -255
rect 164 -261 167 -255
rect 1040 -453 1043 -447
rect 1046 -453 1049 -447
rect 1063 -453 1066 -447
rect 1069 -453 1072 -447
rect 1086 -453 1089 -447
rect 1092 -453 1095 -447
rect 1109 -453 1112 -447
rect 1115 -453 1118 -447
rect 1132 -453 1135 -447
rect 1138 -453 1141 -447
rect 76 -460 79 -454
rect 82 -460 85 -454
rect 99 -460 102 -454
rect 105 -460 108 -454
rect 155 -460 158 -454
rect 161 -460 164 -454
rect 285 -460 288 -454
rect 291 -460 294 -454
rect 308 -460 311 -454
rect 314 -460 317 -454
rect 331 -460 334 -454
rect 337 -460 340 -454
rect 387 -460 390 -454
rect 393 -460 396 -454
rect 531 -460 534 -454
rect 537 -460 540 -454
rect 554 -460 557 -454
rect 560 -460 563 -454
rect 577 -460 580 -454
rect 583 -460 586 -454
rect 600 -460 603 -454
rect 606 -460 609 -454
rect 656 -460 659 -454
rect 662 -460 665 -454
rect 808 -459 811 -453
rect 814 -459 817 -453
rect 831 -459 834 -453
rect 837 -459 840 -453
rect 854 -459 857 -453
rect 860 -459 863 -453
rect 877 -459 880 -453
rect 883 -459 886 -453
rect 900 -459 903 -453
rect 906 -459 909 -453
rect 956 -459 959 -453
rect 962 -459 965 -453
rect 29 -471 32 -465
rect 35 -471 38 -465
rect 220 -470 223 -464
rect 226 -470 229 -464
rect 447 -470 450 -464
rect 453 -470 456 -464
rect 718 -470 721 -464
rect 724 -470 727 -464
<< ndcontact >>
rect 505 458 509 463
rect 519 458 523 463
rect 528 458 532 463
rect 542 458 546 463
rect 551 458 555 463
rect 565 458 569 463
rect 574 458 578 463
rect 588 458 592 463
rect 597 458 601 463
rect 611 458 615 463
rect 30 311 34 316
rect 44 311 48 316
rect 77 312 81 317
rect 91 312 95 317
rect 100 312 104 317
rect 114 312 118 317
rect 156 312 160 317
rect 170 312 174 317
rect 213 312 217 317
rect 227 312 231 317
rect 278 312 282 317
rect 292 312 296 317
rect 301 312 305 317
rect 315 312 319 317
rect 324 312 328 317
rect 338 312 342 317
rect 380 312 384 317
rect 394 312 398 317
rect 441 312 445 317
rect 455 312 459 317
rect 525 312 529 317
rect 539 312 543 317
rect 548 312 552 317
rect 562 312 566 317
rect 571 312 575 317
rect 585 312 589 317
rect 594 312 598 317
rect 608 312 612 317
rect 650 312 654 317
rect 664 312 668 317
rect 715 311 719 316
rect 729 311 733 316
rect 805 312 809 317
rect 819 312 823 317
rect 828 312 832 317
rect 842 312 846 317
rect 851 312 855 317
rect 865 312 869 317
rect 874 312 878 317
rect 888 312 892 317
rect 897 312 901 317
rect 911 312 915 317
rect 953 312 957 317
rect 967 312 971 317
rect 19 152 24 156
rect 33 152 37 156
rect 42 152 47 156
rect 56 152 60 156
rect 73 152 77 156
rect 87 152 91 156
rect 96 152 100 156
rect 110 152 114 156
rect 153 174 157 179
rect 167 174 171 179
rect 18 7 23 11
rect 32 7 36 11
rect 41 7 46 11
rect 55 7 59 11
rect 72 7 76 11
rect 86 7 90 11
rect 95 7 99 11
rect 109 7 113 11
rect 152 29 156 34
rect 166 29 170 34
rect 282 -63 286 -58
rect 296 -63 300 -58
rect 305 -63 309 -58
rect 319 -63 323 -58
rect 328 -63 332 -58
rect 342 -63 346 -58
rect 351 -63 355 -58
rect 365 -63 369 -58
rect 407 -63 411 -58
rect 421 -63 425 -58
rect 18 -155 23 -151
rect 32 -155 36 -151
rect 41 -155 46 -151
rect 55 -155 59 -151
rect 72 -155 76 -151
rect 86 -155 90 -151
rect 95 -155 99 -151
rect 109 -155 113 -151
rect 152 -133 156 -128
rect 166 -133 170 -128
rect 19 -309 24 -305
rect 33 -309 37 -305
rect 42 -309 47 -305
rect 56 -309 60 -305
rect 73 -309 77 -305
rect 87 -309 91 -305
rect 96 -309 100 -305
rect 110 -309 114 -305
rect 153 -287 157 -282
rect 167 -287 171 -282
rect 1035 -481 1039 -476
rect 1049 -481 1053 -476
rect 1058 -481 1062 -476
rect 1072 -481 1076 -476
rect 1081 -481 1085 -476
rect 1095 -481 1099 -476
rect 1104 -481 1108 -476
rect 1118 -481 1122 -476
rect 1127 -481 1131 -476
rect 1141 -481 1145 -476
rect 24 -497 28 -492
rect 38 -497 42 -492
rect 71 -496 75 -491
rect 85 -496 89 -491
rect 94 -496 98 -491
rect 108 -496 112 -491
rect 150 -496 154 -491
rect 164 -496 168 -491
rect 215 -496 219 -491
rect 229 -496 233 -491
rect 280 -496 284 -491
rect 294 -496 298 -491
rect 303 -496 307 -491
rect 317 -496 321 -491
rect 326 -496 330 -491
rect 340 -496 344 -491
rect 382 -496 386 -491
rect 396 -496 400 -491
rect 442 -496 446 -491
rect 456 -496 460 -491
rect 526 -496 530 -491
rect 540 -496 544 -491
rect 549 -496 553 -491
rect 563 -496 567 -491
rect 572 -496 576 -491
rect 586 -496 590 -491
rect 595 -496 599 -491
rect 609 -496 613 -491
rect 651 -496 655 -491
rect 665 -496 669 -491
rect 713 -496 717 -491
rect 727 -496 731 -491
rect 803 -495 807 -490
rect 817 -495 821 -490
rect 826 -495 830 -490
rect 840 -495 844 -490
rect 849 -495 853 -490
rect 863 -495 867 -490
rect 872 -495 876 -490
rect 886 -495 890 -490
rect 895 -495 899 -490
rect 909 -495 913 -490
rect 951 -495 955 -490
rect 965 -495 969 -490
<< pdcontact >>
rect 505 486 510 492
rect 519 486 523 492
rect 528 486 533 492
rect 542 486 546 492
rect 551 486 556 492
rect 565 486 569 492
rect 574 486 579 492
rect 588 486 592 492
rect 597 486 602 492
rect 611 486 615 492
rect 77 348 82 354
rect 91 348 95 354
rect 100 348 105 354
rect 114 348 118 354
rect 156 348 161 354
rect 170 348 174 354
rect 278 348 283 354
rect 292 348 296 354
rect 301 348 306 354
rect 315 348 319 354
rect 324 348 329 354
rect 338 348 342 354
rect 380 348 385 354
rect 394 348 398 354
rect 525 348 530 354
rect 539 348 543 354
rect 548 348 553 354
rect 562 348 566 354
rect 571 348 576 354
rect 585 348 589 354
rect 594 348 599 354
rect 608 348 612 354
rect 650 348 655 354
rect 664 348 668 354
rect 805 348 810 354
rect 819 348 823 354
rect 828 348 833 354
rect 842 348 846 354
rect 851 348 856 354
rect 865 348 869 354
rect 874 348 879 354
rect 888 348 892 354
rect 897 348 902 354
rect 911 348 915 354
rect 953 348 958 354
rect 967 348 971 354
rect 30 337 35 343
rect 44 337 48 343
rect 213 338 218 344
rect 227 338 231 344
rect 441 338 446 344
rect 455 338 459 344
rect 715 337 720 343
rect 729 337 733 343
rect 19 205 24 211
rect 33 205 37 211
rect 42 205 47 211
rect 56 205 60 211
rect 73 205 78 211
rect 87 205 91 211
rect 96 205 101 211
rect 110 205 114 211
rect 153 200 158 206
rect 167 200 171 206
rect 18 60 23 66
rect 32 60 36 66
rect 41 60 46 66
rect 55 60 59 66
rect 72 60 77 66
rect 86 60 90 66
rect 95 60 100 66
rect 109 60 113 66
rect 152 55 157 61
rect 166 55 170 61
rect 282 -27 287 -21
rect 296 -27 300 -21
rect 305 -27 310 -21
rect 319 -27 323 -21
rect 328 -27 333 -21
rect 342 -27 346 -21
rect 351 -27 356 -21
rect 365 -27 369 -21
rect 407 -27 412 -21
rect 421 -27 425 -21
rect 18 -102 23 -96
rect 32 -102 36 -96
rect 41 -102 46 -96
rect 55 -102 59 -96
rect 72 -102 77 -96
rect 86 -102 90 -96
rect 95 -102 100 -96
rect 109 -102 113 -96
rect 152 -107 157 -101
rect 166 -107 170 -101
rect 19 -256 24 -250
rect 33 -256 37 -250
rect 42 -256 47 -250
rect 56 -256 60 -250
rect 73 -256 78 -250
rect 87 -256 91 -250
rect 96 -256 101 -250
rect 110 -256 114 -250
rect 153 -261 158 -255
rect 167 -261 171 -255
rect 1035 -453 1040 -447
rect 1049 -453 1053 -447
rect 1058 -453 1063 -447
rect 1072 -453 1076 -447
rect 1081 -453 1086 -447
rect 1095 -453 1099 -447
rect 1104 -453 1109 -447
rect 1118 -453 1122 -447
rect 1127 -453 1132 -447
rect 1141 -453 1145 -447
rect 71 -460 76 -454
rect 85 -460 89 -454
rect 94 -460 99 -454
rect 108 -460 112 -454
rect 150 -460 155 -454
rect 164 -460 168 -454
rect 280 -460 285 -454
rect 294 -460 298 -454
rect 303 -460 308 -454
rect 317 -460 321 -454
rect 326 -460 331 -454
rect 340 -460 344 -454
rect 382 -460 387 -454
rect 396 -460 400 -454
rect 526 -460 531 -454
rect 540 -460 544 -454
rect 549 -460 554 -454
rect 563 -460 567 -454
rect 572 -460 577 -454
rect 586 -460 590 -454
rect 595 -460 600 -454
rect 609 -460 613 -454
rect 651 -460 656 -454
rect 665 -460 669 -454
rect 803 -459 808 -453
rect 817 -459 821 -453
rect 826 -459 831 -453
rect 840 -459 844 -453
rect 849 -459 854 -453
rect 863 -459 867 -453
rect 872 -459 877 -453
rect 886 -459 890 -453
rect 895 -459 900 -453
rect 909 -459 913 -453
rect 951 -459 956 -453
rect 965 -459 969 -453
rect 24 -471 29 -465
rect 38 -471 42 -465
rect 215 -470 220 -464
rect 229 -470 233 -464
rect 442 -470 447 -464
rect 456 -470 460 -464
rect 713 -470 718 -464
rect 727 -470 731 -464
<< polysilicon >>
rect 513 492 516 496
rect 536 492 539 496
rect 559 492 562 496
rect 582 492 585 496
rect 605 492 608 496
rect 513 463 516 486
rect 536 463 539 486
rect 559 463 562 486
rect 582 463 585 486
rect 605 474 608 486
rect 603 470 608 474
rect 605 463 608 470
rect 513 438 516 458
rect 536 438 539 458
rect 559 438 562 458
rect 582 442 585 458
rect 605 451 608 458
rect 85 354 88 357
rect 108 354 111 357
rect 164 354 167 357
rect 286 354 289 357
rect 309 354 312 357
rect 332 354 335 357
rect 388 354 391 357
rect 533 354 536 357
rect 556 354 559 357
rect 579 354 582 357
rect 602 354 605 357
rect 658 354 661 357
rect 813 354 816 357
rect 836 354 839 357
rect 859 354 862 357
rect 882 354 885 357
rect 905 354 908 357
rect 961 354 964 357
rect 38 343 41 346
rect 38 326 41 337
rect 85 328 88 348
rect 36 322 41 326
rect 83 324 88 328
rect 38 316 41 322
rect 85 317 88 324
rect 108 317 111 348
rect 164 338 167 348
rect 221 344 224 347
rect 286 339 289 348
rect 162 334 167 338
rect 164 317 167 334
rect 221 327 224 338
rect 280 335 289 339
rect 219 323 224 327
rect 221 317 224 323
rect 286 317 289 335
rect 309 333 312 348
rect 307 329 312 333
rect 309 317 312 329
rect 332 328 335 348
rect 388 338 391 348
rect 449 344 452 347
rect 533 339 536 348
rect 386 334 391 338
rect 330 324 335 328
rect 332 317 335 324
rect 388 317 391 334
rect 449 327 452 338
rect 530 335 536 339
rect 447 323 452 327
rect 449 317 452 323
rect 533 317 536 335
rect 556 333 559 348
rect 554 329 559 333
rect 556 317 559 329
rect 579 325 582 348
rect 577 321 582 325
rect 579 317 582 321
rect 602 317 605 348
rect 658 338 661 348
rect 723 343 726 346
rect 656 334 661 338
rect 658 317 661 334
rect 723 326 726 337
rect 813 328 816 348
rect 721 322 726 326
rect 811 324 816 328
rect 723 316 726 322
rect 813 317 816 324
rect 836 317 839 348
rect 859 317 862 348
rect 882 317 885 348
rect 905 317 908 348
rect 961 338 964 348
rect 959 334 964 338
rect 961 317 964 334
rect 38 304 41 311
rect 85 308 88 312
rect 108 296 111 312
rect 164 308 167 312
rect 221 305 224 312
rect 286 308 289 312
rect 309 308 312 312
rect 332 308 335 312
rect 388 308 391 312
rect 449 305 452 312
rect 533 308 536 312
rect 556 308 559 312
rect 579 308 582 312
rect 85 293 111 296
rect 602 293 605 312
rect 658 308 661 312
rect 723 304 726 311
rect 813 308 816 312
rect 3 230 53 233
rect 3 135 6 230
rect 27 211 30 215
rect 50 211 53 230
rect 81 211 84 292
rect 836 284 839 312
rect 859 284 862 312
rect 882 283 885 312
rect 905 284 908 312
rect 961 308 964 312
rect 104 211 107 250
rect 161 206 164 209
rect 27 166 30 205
rect 50 199 53 205
rect 81 187 84 205
rect 104 187 107 205
rect 161 189 164 200
rect 79 183 84 187
rect 97 183 107 187
rect 27 163 53 166
rect 27 156 30 160
rect 50 156 53 163
rect 81 156 84 183
rect 104 156 107 183
rect 159 185 164 189
rect 27 135 30 152
rect 50 148 53 152
rect 81 149 84 152
rect 104 150 107 152
rect 92 148 107 150
rect 50 146 72 148
rect 70 144 72 146
rect 92 144 94 148
rect 70 142 94 144
rect 123 135 126 183
rect 161 179 164 185
rect 161 167 164 174
rect 3 132 126 135
rect 93 118 96 121
rect -61 115 96 118
rect -61 114 83 115
rect 2 85 52 88
rect 2 -10 5 85
rect 26 66 29 70
rect 49 66 52 85
rect 80 66 83 114
rect 103 66 106 112
rect 160 61 163 64
rect 26 42 29 60
rect 49 54 52 60
rect 80 42 83 60
rect 103 42 106 60
rect 160 44 163 55
rect 15 38 29 42
rect 78 38 83 42
rect 96 38 106 42
rect 26 21 29 38
rect 26 18 52 21
rect 26 11 29 15
rect 49 11 52 18
rect 80 11 83 38
rect 103 11 106 38
rect 158 40 163 44
rect 26 -10 29 7
rect 49 3 52 7
rect 80 4 83 7
rect 103 5 106 7
rect 91 3 106 5
rect 49 1 71 3
rect 69 -1 71 1
rect 91 -1 93 3
rect 69 -3 93 -1
rect 122 -10 125 38
rect 160 34 163 40
rect 160 22 163 29
rect 2 -13 125 -10
rect 290 -21 293 -18
rect 313 -21 316 -18
rect 336 -21 339 -18
rect 359 -21 362 -18
rect 415 -21 418 -18
rect -90 -47 83 -44
rect 80 -50 83 -47
rect 2 -77 52 -74
rect 2 -172 5 -77
rect 26 -96 29 -92
rect 49 -96 52 -77
rect 80 -96 83 -55
rect 103 -96 106 -31
rect 290 -47 293 -27
rect 288 -51 293 -47
rect 290 -58 293 -51
rect 313 -58 316 -27
rect 336 -58 339 -27
rect 359 -58 362 -27
rect 415 -37 418 -27
rect 413 -41 418 -37
rect 415 -58 418 -41
rect 290 -67 293 -63
rect 313 -78 316 -63
rect 336 -78 339 -63
rect 359 -79 362 -63
rect 415 -67 418 -63
rect 160 -101 163 -98
rect 26 -119 29 -102
rect 49 -108 52 -102
rect 15 -123 29 -119
rect 80 -120 83 -102
rect 103 -120 106 -102
rect 160 -118 163 -107
rect 26 -141 29 -123
rect 78 -124 83 -120
rect 96 -124 106 -120
rect 26 -144 52 -141
rect 26 -151 29 -147
rect 49 -151 52 -144
rect 80 -151 83 -124
rect 103 -151 106 -124
rect 158 -122 163 -118
rect 26 -172 29 -155
rect 49 -159 52 -155
rect 80 -158 83 -155
rect 103 -157 106 -155
rect 91 -159 106 -157
rect 49 -161 71 -159
rect 69 -163 71 -161
rect 91 -163 93 -159
rect 69 -165 93 -163
rect 122 -172 125 -124
rect 160 -128 163 -122
rect 160 -140 163 -133
rect 2 -175 125 -172
rect -118 -199 81 -196
rect 3 -231 53 -228
rect 3 -326 6 -231
rect 27 -250 30 -246
rect 50 -250 53 -231
rect 81 -250 84 -199
rect 104 -250 107 -209
rect 161 -255 164 -252
rect 27 -295 30 -256
rect 50 -262 53 -256
rect 81 -274 84 -256
rect 104 -274 107 -256
rect 161 -272 164 -261
rect 79 -278 84 -274
rect 97 -278 107 -274
rect 27 -298 53 -295
rect 27 -305 30 -301
rect 50 -305 53 -298
rect 81 -305 84 -278
rect 104 -305 107 -278
rect 159 -276 164 -272
rect 27 -326 30 -309
rect 50 -313 53 -309
rect 81 -312 84 -309
rect 104 -311 107 -309
rect 92 -313 107 -311
rect 50 -315 72 -313
rect 70 -317 72 -315
rect 92 -317 94 -313
rect 70 -319 94 -317
rect 123 -326 126 -278
rect 161 -282 164 -276
rect 161 -294 164 -287
rect 3 -329 126 -326
rect 79 -454 82 -451
rect 102 -454 105 -451
rect 158 -454 161 -451
rect 288 -454 291 -451
rect 311 -454 314 -451
rect 334 -454 337 -373
rect 580 -392 583 -373
rect 580 -396 633 -392
rect 390 -454 393 -451
rect 534 -454 537 -451
rect 557 -454 560 -451
rect 580 -454 583 -396
rect 603 -454 606 -427
rect 659 -454 662 -451
rect 811 -453 814 -450
rect 834 -453 837 -418
rect 857 -453 860 -440
rect 880 -453 883 -439
rect 903 -453 906 -438
rect 1043 -447 1046 -443
rect 1066 -447 1069 -443
rect 1089 -447 1092 -443
rect 1112 -447 1115 -443
rect 1135 -447 1138 -443
rect 959 -453 962 -450
rect 32 -465 35 -462
rect 32 -482 35 -471
rect 79 -480 82 -460
rect 30 -486 35 -482
rect 77 -484 82 -480
rect 32 -492 35 -486
rect 79 -491 82 -484
rect 102 -491 105 -460
rect 158 -470 161 -460
rect 223 -464 226 -461
rect 288 -469 291 -460
rect 156 -474 161 -470
rect 158 -491 161 -474
rect 223 -481 226 -470
rect 282 -473 291 -469
rect 221 -485 226 -481
rect 223 -491 226 -485
rect 288 -491 291 -473
rect 311 -475 314 -460
rect 309 -479 314 -475
rect 311 -491 314 -479
rect 334 -491 337 -460
rect 390 -470 393 -460
rect 450 -464 453 -461
rect 534 -469 537 -460
rect 388 -474 393 -470
rect 390 -491 393 -474
rect 450 -481 453 -470
rect 531 -473 537 -469
rect 448 -485 453 -481
rect 450 -491 453 -485
rect 534 -491 537 -473
rect 557 -491 560 -460
rect 580 -491 583 -460
rect 603 -491 606 -460
rect 659 -470 662 -460
rect 721 -464 724 -461
rect 657 -474 662 -470
rect 659 -491 662 -474
rect 721 -481 724 -470
rect 811 -479 814 -459
rect 719 -485 724 -481
rect 809 -483 814 -479
rect 721 -491 724 -485
rect 811 -490 814 -483
rect 834 -490 837 -459
rect 857 -490 860 -459
rect 880 -490 883 -459
rect 903 -490 906 -459
rect 959 -469 962 -459
rect 1043 -467 1046 -453
rect 957 -473 962 -469
rect 1035 -471 1046 -467
rect 959 -490 962 -473
rect 1043 -476 1046 -471
rect 1066 -476 1069 -453
rect 1089 -476 1092 -453
rect 1112 -476 1115 -453
rect 1135 -465 1138 -453
rect 1133 -469 1138 -465
rect 1135 -476 1138 -469
rect 1043 -485 1046 -481
rect 32 -504 35 -497
rect 79 -500 82 -496
rect 102 -532 105 -496
rect 158 -500 161 -496
rect 223 -503 226 -496
rect 288 -500 291 -496
rect 311 -500 314 -496
rect 334 -500 337 -496
rect 390 -500 393 -496
rect 450 -503 453 -496
rect 534 -500 537 -496
rect 557 -521 560 -496
rect 580 -500 583 -496
rect 603 -500 606 -496
rect 659 -500 662 -496
rect 721 -503 724 -496
rect 811 -499 814 -495
rect 834 -501 837 -495
rect 857 -501 860 -495
rect 880 -501 883 -495
rect 903 -501 906 -495
rect 959 -499 962 -495
rect 1066 -501 1069 -481
rect 1089 -501 1092 -481
rect 1112 -497 1115 -481
rect 1135 -488 1138 -481
<< polycontact >>
rect 598 470 603 474
rect 512 433 516 438
rect 535 433 539 438
rect 559 433 563 438
rect 582 437 586 442
rect 31 322 36 326
rect 78 324 83 328
rect 157 334 162 338
rect 275 335 280 339
rect 214 323 219 327
rect 302 329 307 333
rect 381 334 386 338
rect 325 324 330 328
rect 525 335 530 339
rect 442 323 447 327
rect 549 329 554 333
rect 572 321 577 325
rect 651 334 656 338
rect 716 322 721 326
rect 806 324 811 328
rect 954 334 959 338
rect 80 292 85 296
rect 601 289 606 293
rect 834 278 839 284
rect 858 278 863 284
rect 880 277 885 283
rect 904 278 909 284
rect 103 250 108 254
rect 74 183 79 187
rect 123 183 127 188
rect 154 185 159 189
rect 93 121 98 125
rect -66 114 -61 118
rect 103 112 108 116
rect 10 38 15 42
rect 73 38 78 42
rect 122 38 126 43
rect 153 40 158 44
rect 103 -31 107 -26
rect -94 -47 -90 -42
rect 80 -55 84 -50
rect 283 -51 288 -47
rect 408 -41 413 -37
rect 312 -82 317 -78
rect 335 -82 340 -78
rect 358 -83 363 -79
rect 10 -123 15 -119
rect 73 -124 78 -120
rect 122 -124 126 -119
rect 153 -122 158 -118
rect -123 -199 -118 -195
rect 81 -199 86 -195
rect 103 -209 108 -205
rect 74 -278 79 -274
rect 123 -278 127 -273
rect 154 -276 159 -272
rect 333 -373 338 -369
rect 578 -373 583 -369
rect 633 -396 638 -392
rect 831 -418 837 -414
rect 600 -427 606 -423
rect 855 -440 861 -436
rect 879 -439 885 -435
rect 901 -438 907 -434
rect 25 -486 30 -482
rect 72 -484 77 -480
rect 151 -474 156 -470
rect 277 -473 282 -469
rect 216 -485 221 -481
rect 304 -479 309 -475
rect 383 -474 388 -470
rect 526 -473 531 -469
rect 443 -485 448 -481
rect 652 -474 657 -470
rect 714 -485 719 -481
rect 804 -483 809 -479
rect 952 -473 957 -469
rect 1029 -472 1035 -467
rect 1128 -469 1133 -465
rect 1065 -506 1069 -501
rect 1089 -506 1093 -501
rect 1112 -502 1116 -497
rect 557 -525 562 -521
rect 101 -537 107 -532
<< metal1 >>
rect -12 500 602 504
rect -12 499 510 500
rect -33 304 -28 447
rect -12 364 -7 499
rect 505 492 510 499
rect 597 492 602 500
rect 523 486 528 492
rect 546 486 551 492
rect 569 486 574 492
rect 588 474 592 486
rect 611 474 615 486
rect 519 470 598 474
rect 611 470 621 474
rect 519 463 523 470
rect 542 463 546 470
rect 565 463 569 470
rect 588 463 592 470
rect 611 463 615 470
rect 505 451 509 458
rect 528 451 532 458
rect 551 451 555 458
rect 574 451 578 458
rect 597 451 601 458
rect 41 447 601 451
rect 642 446 985 450
rect 182 433 512 438
rect 182 376 186 433
rect 535 425 539 433
rect 642 441 646 446
rect 586 437 646 441
rect 559 429 681 433
rect 406 422 539 425
rect 406 375 409 422
rect 678 372 681 429
rect -12 361 977 364
rect -12 360 404 361
rect -33 299 -32 304
rect -50 270 -45 271
rect -123 -611 -119 -199
rect -110 -603 -106 -124
rect -94 -588 -90 -47
rect -78 -563 -73 37
rect -66 -547 -61 114
rect -50 -532 -45 265
rect -42 -518 -37 291
rect -33 125 -28 299
rect -12 257 -7 360
rect 23 354 27 360
rect 77 354 82 360
rect 100 354 105 360
rect 156 354 161 360
rect 206 355 211 360
rect 23 349 54 354
rect 30 343 35 349
rect 206 350 237 355
rect 278 354 283 360
rect 301 354 306 360
rect 324 354 329 360
rect 380 354 385 360
rect 434 355 439 361
rect 495 360 977 361
rect 44 326 48 337
rect 91 338 95 348
rect 114 338 118 348
rect 170 338 174 348
rect 213 344 218 350
rect 434 350 465 355
rect 525 354 530 360
rect 548 354 553 360
rect 571 354 576 360
rect 594 354 599 360
rect 650 354 655 360
rect 708 354 712 360
rect 805 354 810 360
rect 828 354 833 360
rect 851 354 856 360
rect 874 354 879 360
rect 897 354 902 360
rect 953 354 958 360
rect 91 334 157 338
rect 170 334 180 338
rect 292 339 296 348
rect 315 339 319 348
rect 338 339 342 348
rect 53 326 78 328
rect 1 322 31 326
rect 44 324 78 326
rect 44 322 57 324
rect 1 270 5 322
rect 44 316 48 322
rect 114 317 118 334
rect 170 317 174 334
rect 227 327 231 338
rect 238 335 275 339
rect 292 338 342 339
rect 394 338 398 348
rect 441 344 446 350
rect 708 349 739 354
rect 292 336 381 338
rect 238 327 241 335
rect 338 334 381 336
rect 394 334 404 338
rect 539 339 543 348
rect 562 339 566 348
rect 585 339 589 348
rect 608 339 612 348
rect 186 323 214 327
rect 227 323 241 327
rect 244 329 302 332
rect 227 317 231 323
rect 244 320 247 329
rect 322 326 325 327
rect 95 312 100 317
rect 236 317 247 320
rect 256 323 325 326
rect 236 312 239 317
rect 30 303 34 311
rect 77 303 81 312
rect 156 303 160 312
rect 213 303 217 312
rect 256 311 259 323
rect 338 317 342 334
rect 394 317 398 334
rect 455 327 459 338
rect 468 335 525 339
rect 539 338 612 339
rect 664 338 668 348
rect 715 343 720 349
rect 539 336 651 338
rect 468 327 472 335
rect 608 334 651 336
rect 664 334 677 338
rect 413 323 442 327
rect 455 323 472 327
rect 475 329 549 332
rect 455 317 459 323
rect 475 319 478 329
rect 250 308 259 311
rect 296 312 301 317
rect 319 312 324 317
rect 464 316 478 319
rect 483 321 572 325
rect 278 303 282 312
rect 380 303 384 312
rect 441 303 445 312
rect 464 311 468 316
rect 483 311 486 321
rect 608 317 612 334
rect 664 317 668 334
rect 729 326 733 337
rect 819 338 823 348
rect 842 338 846 348
rect 865 338 869 348
rect 888 338 892 348
rect 911 338 915 348
rect 967 338 971 348
rect 981 338 985 446
rect 819 334 954 338
rect 967 334 985 338
rect 796 326 806 328
rect 701 322 716 326
rect 729 323 806 326
rect 729 322 797 323
rect 543 312 548 317
rect 566 312 571 317
rect 589 312 594 317
rect 729 316 733 322
rect 911 317 915 334
rect 967 317 971 334
rect 525 303 529 312
rect 650 303 654 312
rect 823 312 828 317
rect 846 312 851 317
rect 869 312 874 317
rect 892 312 897 317
rect 715 303 719 311
rect 805 303 809 312
rect 953 303 957 312
rect 27 300 957 303
rect 654 299 806 300
rect 47 293 80 296
rect 602 276 605 289
rect 1 263 6 265
rect 215 269 407 274
rect 515 271 605 276
rect 1 260 107 263
rect 104 254 107 260
rect 215 262 219 269
rect -33 -24 -29 120
rect -12 112 -8 252
rect 60 244 138 247
rect 19 236 68 240
rect 19 211 24 236
rect 19 156 24 205
rect 33 221 55 226
rect 33 211 37 221
rect 56 211 60 221
rect 33 156 37 205
rect 42 156 47 205
rect 56 156 60 205
rect 65 187 68 236
rect 78 223 96 228
rect 73 211 78 223
rect 96 211 101 223
rect 65 183 74 187
rect 87 178 91 205
rect 65 174 91 178
rect 42 144 47 152
rect 65 144 68 174
rect 87 156 91 174
rect 110 188 114 205
rect 134 189 138 244
rect 151 212 177 217
rect 153 206 158 212
rect 167 189 171 200
rect 110 183 123 188
rect 134 185 154 189
rect 167 185 201 189
rect 110 156 114 183
rect 167 179 171 185
rect 153 166 157 174
rect 42 141 68 144
rect 145 163 177 166
rect 73 141 77 152
rect 96 141 100 152
rect 73 140 100 141
rect 145 140 148 163
rect 73 137 148 140
rect 84 124 88 137
rect 11 121 88 124
rect 98 122 190 125
rect 108 112 180 116
rect -33 -186 -29 -29
rect -12 -37 -8 107
rect 59 99 137 102
rect 18 91 67 95
rect 18 66 23 91
rect 0 38 10 41
rect 18 11 23 60
rect 32 76 54 81
rect 32 66 36 76
rect 55 66 59 76
rect 32 11 36 60
rect 41 11 46 60
rect 55 11 59 60
rect 64 42 67 91
rect 77 78 95 83
rect 72 66 77 78
rect 95 66 100 78
rect 64 38 73 42
rect 86 33 90 60
rect 64 29 90 33
rect 41 -1 46 7
rect 64 -1 67 29
rect 86 11 90 29
rect 109 43 113 60
rect 133 44 137 99
rect 150 67 176 72
rect 152 61 157 67
rect 166 44 170 55
rect 109 38 122 43
rect 133 40 153 44
rect 166 40 187 44
rect 109 11 113 38
rect 166 34 170 40
rect 152 21 156 29
rect 41 -4 67 -1
rect 144 18 176 21
rect 72 -4 76 7
rect 95 -4 99 7
rect 72 -5 99 -4
rect 144 -5 147 18
rect 72 -8 147 -5
rect 83 -24 87 -8
rect 11 -27 87 -24
rect 107 -30 144 -27
rect 169 -37 174 -15
rect -12 -41 174 -37
rect -12 -50 -8 -41
rect 84 -54 163 -51
rect -33 -338 -29 -191
rect -12 -204 -8 -55
rect 59 -63 137 -60
rect 18 -71 67 -67
rect 18 -96 23 -71
rect 0 -123 10 -120
rect 18 -151 23 -102
rect 32 -86 54 -81
rect 32 -96 36 -86
rect 55 -96 59 -86
rect 32 -151 36 -102
rect 41 -151 46 -102
rect 55 -151 59 -102
rect 64 -120 67 -71
rect 77 -84 95 -79
rect 72 -96 77 -84
rect 95 -96 100 -84
rect 64 -124 73 -120
rect 86 -129 90 -102
rect 64 -133 90 -129
rect 41 -163 46 -155
rect 64 -163 67 -133
rect 86 -151 90 -133
rect 109 -119 113 -102
rect 133 -118 137 -63
rect 150 -95 176 -90
rect 152 -101 157 -95
rect 187 -100 192 40
rect 202 -47 208 185
rect 215 -25 218 262
rect 460 258 465 269
rect 227 252 465 258
rect 227 -23 231 252
rect 482 243 485 269
rect 239 238 482 242
rect 239 190 243 238
rect 244 185 435 190
rect 515 176 520 271
rect 515 175 650 176
rect 241 169 650 175
rect 242 45 247 169
rect 695 147 701 278
rect 452 141 701 147
rect 722 278 834 284
rect 247 40 431 45
rect 280 -15 431 -11
rect 282 -21 287 -15
rect 305 -21 310 -15
rect 328 -21 333 -15
rect 351 -21 356 -15
rect 407 -21 412 -15
rect 296 -37 300 -27
rect 319 -37 323 -27
rect 342 -37 346 -27
rect 365 -37 369 -27
rect 421 -37 425 -27
rect 296 -41 408 -37
rect 421 -41 431 -37
rect 202 -51 283 -47
rect 365 -58 369 -41
rect 421 -58 425 -41
rect 277 -63 282 -58
rect 300 -63 305 -58
rect 323 -63 328 -58
rect 346 -63 351 -58
rect 277 -70 281 -63
rect 407 -72 411 -63
rect 281 -75 411 -72
rect 312 -100 317 -82
rect 187 -106 317 -100
rect 166 -118 170 -107
rect 336 -117 340 -82
rect 179 -118 336 -117
rect 109 -124 122 -119
rect 133 -122 153 -118
rect 166 -122 336 -118
rect 359 -120 363 -83
rect 109 -151 113 -124
rect 166 -128 170 -122
rect 152 -141 156 -133
rect 41 -166 67 -163
rect 144 -144 176 -141
rect 72 -166 76 -155
rect 95 -166 99 -155
rect 72 -167 99 -166
rect 144 -167 147 -144
rect 72 -170 147 -167
rect 83 -184 87 -170
rect 83 -186 275 -184
rect 11 -189 275 -186
rect 86 -198 297 -195
rect 108 -209 298 -206
rect -33 -505 -29 -343
rect -12 -444 -8 -209
rect 60 -217 138 -214
rect 19 -225 68 -221
rect 19 -250 24 -225
rect 19 -305 24 -256
rect 33 -240 55 -235
rect 33 -250 37 -240
rect 56 -250 60 -240
rect 33 -305 37 -256
rect 42 -305 47 -256
rect 56 -305 60 -256
rect 65 -274 68 -225
rect 78 -238 96 -233
rect 73 -250 78 -238
rect 96 -250 101 -238
rect 65 -278 74 -274
rect 87 -283 91 -256
rect 65 -287 91 -283
rect 42 -317 47 -309
rect 65 -317 68 -287
rect 87 -305 91 -287
rect 110 -273 114 -256
rect 134 -272 138 -217
rect 151 -249 177 -244
rect 153 -255 158 -249
rect 167 -272 171 -261
rect 359 -271 364 -120
rect 452 -204 456 141
rect 722 130 729 278
rect 858 243 861 278
rect 740 239 861 243
rect 880 176 885 277
rect 744 169 885 176
rect 903 278 904 283
rect 465 126 729 130
rect 465 -193 469 126
rect 903 106 909 278
rect 478 100 909 106
rect 478 99 907 100
rect 478 -117 483 99
rect 532 75 533 79
rect 180 -272 365 -271
rect 110 -278 123 -273
rect 134 -276 154 -272
rect 167 -276 365 -272
rect 110 -305 114 -278
rect 167 -282 171 -276
rect 323 -277 365 -276
rect 153 -295 157 -287
rect 42 -320 68 -317
rect 145 -298 177 -295
rect 73 -320 77 -309
rect 96 -320 100 -309
rect 73 -321 100 -320
rect 145 -321 148 -298
rect 73 -324 148 -321
rect 85 -340 89 -324
rect 11 -343 89 -340
rect 532 -369 540 75
rect 596 45 602 46
rect 560 40 604 45
rect 338 -370 543 -369
rect 338 -373 578 -370
rect 598 -423 604 40
rect 619 -414 623 -210
rect 650 -370 656 -122
rect 650 -376 906 -370
rect 638 -396 884 -392
rect 619 -418 831 -414
rect 598 -427 600 -423
rect 606 -427 860 -423
rect 856 -436 860 -427
rect 879 -435 884 -396
rect 901 -434 906 -376
rect 1003 -439 1132 -435
rect 1003 -440 1040 -439
rect 1003 -443 1008 -440
rect 688 -444 1008 -443
rect -12 -447 1008 -444
rect 1035 -447 1040 -440
rect 1127 -447 1132 -439
rect -12 -448 406 -447
rect 17 -454 21 -448
rect 71 -454 76 -448
rect 94 -454 99 -448
rect 150 -454 155 -448
rect 208 -453 213 -448
rect 17 -459 48 -454
rect 24 -465 29 -459
rect 208 -458 239 -453
rect 280 -454 285 -448
rect 303 -454 308 -448
rect 326 -454 331 -448
rect 382 -454 387 -448
rect 435 -453 440 -447
rect 496 -448 692 -447
rect 38 -482 42 -471
rect 85 -470 89 -460
rect 108 -470 112 -460
rect 164 -470 168 -460
rect 215 -464 220 -458
rect 435 -458 466 -453
rect 526 -454 531 -448
rect 549 -454 554 -448
rect 572 -454 577 -448
rect 595 -454 600 -448
rect 651 -454 656 -448
rect 706 -453 710 -447
rect 803 -453 808 -447
rect 826 -453 831 -447
rect 849 -453 854 -447
rect 872 -453 877 -447
rect 895 -453 900 -447
rect 951 -453 956 -447
rect 1053 -453 1058 -447
rect 1076 -453 1081 -447
rect 1099 -453 1104 -447
rect 85 -474 151 -470
rect 164 -474 172 -470
rect 294 -469 298 -460
rect 317 -469 321 -460
rect 340 -469 344 -460
rect 47 -482 72 -480
rect 8 -486 25 -482
rect 38 -484 72 -482
rect 38 -486 51 -484
rect 38 -492 42 -486
rect 108 -491 112 -474
rect 164 -491 168 -474
rect 229 -481 233 -470
rect 240 -473 277 -469
rect 294 -470 344 -469
rect 396 -470 400 -460
rect 442 -464 447 -458
rect 706 -458 737 -453
rect 294 -472 383 -470
rect 240 -481 243 -473
rect 340 -474 383 -472
rect 396 -474 403 -470
rect 540 -469 544 -460
rect 563 -469 567 -460
rect 586 -469 590 -460
rect 609 -469 613 -460
rect 199 -485 216 -481
rect 229 -485 243 -481
rect 246 -479 304 -476
rect 229 -491 233 -485
rect 246 -488 249 -479
rect 89 -496 94 -491
rect 238 -491 249 -488
rect 340 -491 344 -474
rect 396 -491 400 -474
rect 456 -481 460 -470
rect 469 -473 526 -469
rect 540 -470 613 -469
rect 665 -470 669 -460
rect 713 -464 718 -458
rect 540 -472 652 -470
rect 469 -481 473 -473
rect 419 -485 443 -481
rect 456 -485 473 -481
rect 609 -474 652 -472
rect 665 -474 678 -470
rect 456 -491 460 -485
rect 609 -491 613 -474
rect 665 -491 669 -474
rect 727 -481 731 -470
rect 817 -469 821 -459
rect 840 -469 844 -459
rect 863 -469 867 -459
rect 886 -469 890 -459
rect 909 -469 913 -459
rect 965 -468 969 -459
rect 1118 -465 1122 -453
rect 1141 -465 1145 -453
rect 817 -473 952 -469
rect 965 -472 1029 -468
rect 1049 -469 1128 -465
rect 1141 -469 1151 -465
rect 794 -481 804 -479
rect 699 -485 714 -481
rect 727 -484 804 -481
rect 727 -485 795 -484
rect 727 -491 731 -485
rect 909 -490 913 -473
rect 965 -490 969 -472
rect 1049 -476 1053 -469
rect 1072 -476 1076 -469
rect 1095 -476 1099 -469
rect 1118 -476 1122 -469
rect 1141 -476 1145 -469
rect 1035 -488 1039 -481
rect 1058 -488 1062 -481
rect 1081 -488 1085 -481
rect 1104 -488 1108 -481
rect 1127 -488 1131 -481
rect 238 -496 241 -491
rect 298 -496 303 -491
rect 321 -496 326 -491
rect 544 -496 549 -491
rect 567 -496 572 -491
rect 590 -496 595 -491
rect 821 -495 826 -490
rect 844 -495 849 -490
rect 867 -495 872 -490
rect 890 -495 895 -490
rect 1026 -492 1131 -488
rect 24 -505 28 -497
rect 71 -505 75 -496
rect 150 -505 154 -496
rect 215 -505 219 -496
rect 280 -505 284 -496
rect 382 -505 386 -496
rect 442 -505 446 -496
rect 526 -505 530 -496
rect 651 -505 655 -496
rect 713 -504 717 -496
rect 803 -504 807 -495
rect 951 -503 955 -495
rect 1026 -503 1030 -492
rect 951 -504 1030 -503
rect 688 -505 1030 -504
rect -33 -507 1030 -505
rect -33 -508 804 -507
rect -42 -523 2 -518
rect -50 -537 101 -532
rect 193 -547 198 -521
rect -66 -552 198 -547
rect 236 -563 241 -520
rect -78 -569 241 -563
rect 414 -588 419 -526
rect -94 -593 419 -588
rect 700 -525 701 -523
rect 557 -601 561 -525
rect 534 -602 561 -601
rect 348 -603 561 -602
rect -110 -606 561 -603
rect 696 -611 701 -525
rect 1065 -529 1069 -506
rect 719 -534 1069 -529
rect 1089 -540 1093 -506
rect 720 -545 1093 -540
rect 1089 -546 1093 -545
rect 1112 -570 1116 -502
rect 726 -575 1116 -570
rect -123 -615 701 -611
<< m2contact >>
rect -33 447 -28 452
rect 36 447 41 452
rect 181 371 186 376
rect 405 370 410 375
rect 677 367 682 372
rect -32 299 -27 304
rect -42 291 -37 296
rect -50 265 -45 270
rect -78 37 -73 42
rect -110 -124 -105 -119
rect -33 120 -28 125
rect 180 334 185 339
rect 404 334 409 339
rect 181 322 186 327
rect 22 299 27 304
rect 235 307 240 312
rect 245 307 250 312
rect 677 334 682 339
rect 408 322 413 327
rect 695 321 701 326
rect 464 306 469 311
rect 481 306 486 311
rect 42 292 47 297
rect 1 265 6 270
rect 407 269 412 274
rect 460 269 465 274
rect 481 269 486 274
rect 695 278 701 283
rect -12 252 -7 257
rect 55 243 60 248
rect 55 221 60 226
rect 73 223 78 228
rect 96 223 101 228
rect 146 212 151 217
rect 201 185 208 190
rect 6 120 11 125
rect 190 122 195 127
rect -12 107 -7 112
rect 180 111 185 116
rect -33 -29 -28 -24
rect 54 98 59 103
rect -5 37 0 42
rect 54 76 59 81
rect 72 78 77 83
rect 95 78 100 83
rect 145 67 150 72
rect 187 40 192 45
rect 6 -29 11 -24
rect 169 -15 174 -10
rect 144 -30 149 -25
rect -12 -55 -7 -50
rect 163 -55 168 -50
rect -33 -191 -28 -186
rect 54 -64 59 -59
rect -5 -124 0 -119
rect 54 -86 59 -81
rect 72 -84 77 -79
rect 95 -84 100 -79
rect 145 -95 150 -90
rect 482 238 487 243
rect 237 185 244 190
rect 435 185 440 190
rect 650 169 659 176
rect 242 40 247 45
rect 431 40 436 45
rect 275 -15 280 -10
rect 214 -30 219 -25
rect 227 -28 232 -23
rect 276 -75 281 -70
rect 336 -122 341 -117
rect 6 -191 11 -186
rect 275 -189 280 -184
rect 297 -198 302 -193
rect -12 -209 -7 -204
rect 298 -209 303 -204
rect -33 -343 -28 -338
rect 55 -218 60 -213
rect 55 -240 60 -235
rect 73 -238 78 -233
rect 96 -238 101 -233
rect 146 -249 151 -244
rect 734 239 740 244
rect 739 169 744 176
rect 478 -122 483 -117
rect 533 75 542 82
rect 464 -198 469 -193
rect 451 -209 456 -204
rect 6 -343 11 -338
rect 554 40 560 45
rect 649 -122 657 -117
rect 619 -210 624 -205
rect 172 -474 178 -469
rect 3 -487 8 -482
rect 403 -474 408 -469
rect 193 -486 199 -481
rect 414 -485 419 -480
rect 678 -474 683 -469
rect 693 -486 699 -481
rect 237 -501 242 -496
rect 2 -523 7 -518
rect 193 -521 198 -516
rect 236 -520 241 -515
rect 414 -526 419 -521
rect 694 -525 700 -520
rect 713 -534 719 -529
rect 714 -545 720 -540
rect 720 -575 726 -570
<< metal2 >>
rect -28 448 36 451
rect 181 339 184 371
rect 405 339 408 370
rect 678 339 681 367
rect -27 300 22 303
rect -37 292 42 295
rect -45 266 1 270
rect -7 252 77 257
rect 56 226 59 243
rect 73 228 77 252
rect 101 224 150 227
rect 147 217 150 224
rect -28 120 6 124
rect 181 116 185 322
rect 235 295 238 307
rect 190 292 238 295
rect 190 127 194 292
rect 245 286 249 307
rect 202 280 249 286
rect 202 190 208 280
rect 408 274 411 322
rect 460 274 464 309
rect 481 274 485 306
rect 696 283 699 321
rect 487 239 734 243
rect 208 185 237 189
rect 440 185 539 190
rect -7 107 77 112
rect 55 81 58 98
rect 73 83 77 107
rect 533 82 539 185
rect 659 169 739 176
rect 100 79 149 82
rect 146 72 149 79
rect -73 38 -5 41
rect 192 40 242 45
rect 436 40 554 45
rect 174 -14 275 -10
rect -28 -29 6 -25
rect 149 -30 214 -27
rect -7 -55 76 -50
rect 227 -51 232 -28
rect 168 -54 232 -51
rect 55 -81 58 -64
rect 72 -79 76 -55
rect 100 -83 149 -80
rect 146 -90 149 -83
rect -105 -124 -5 -120
rect 276 -184 280 -75
rect 341 -122 478 -117
rect 483 -122 649 -117
rect -28 -191 6 -187
rect 302 -198 464 -194
rect -7 -209 78 -204
rect 303 -209 451 -205
rect 456 -209 619 -205
rect 56 -235 59 -218
rect 74 -233 78 -209
rect 101 -237 150 -234
rect 147 -244 150 -237
rect -28 -343 6 -339
rect 3 -518 7 -487
rect 173 -571 176 -474
rect 193 -516 198 -486
rect 237 -515 240 -501
rect 404 -536 407 -474
rect 414 -521 418 -485
rect 679 -530 682 -474
rect 694 -520 697 -486
rect 679 -534 713 -530
rect 404 -539 602 -536
rect 598 -542 602 -539
rect 598 -545 714 -542
rect 173 -575 720 -571
<< labels >>
rlabel metal1 84 137 89 139 1 gnd
rlabel metal1 90 224 93 227 1 vdd
rlabel polysilicon 80 184 83 187 1 A3
rlabel polysilicon 101 184 104 187 1 B3
rlabel polysilicon 79 38 82 41 1 A2
rlabel polysilicon 99 39 102 42 1 B2
rlabel polysilicon 79 -123 82 -120 1 A1
rlabel polysilicon 99 -123 102 -120 1 B1
rlabel polysilicon 80 -277 83 -274 1 A0
rlabel polysilicon 99 -277 102 -274 1 B0
rlabel metal1 617 471 620 473 1 AB
rlabel metal1 427 -40 430 -38 1 AequalB
rlabel metal1 1147 -468 1150 -466 7 BA
<< end >>
